module TEMAC_CORE_aead6cd6dadd(reset, mac_has_sgmii, rx_correct_frame, rx_error_frame, rx_data, rx_data_vld, rx_status_vector, rx_status_vld, rx_clk_en, tx_data, tx_data_en, tx_stop, tx_rdy, tx_retransmit, tx_collision, tx_clk_en, tx_ifg_val, tx_status_vector, tx_status_vld, pause_req, pause_val,
tx_mac_clk, rx_mac_clk, speed_1000,speed_100, speed_10, gmii_col, gmii_crs, gmii_tx_clken, gmii_txd, gmii_tx_en, gmii_tx_er, gmii_rxd, gmii_rx_vld, gmii_rx_er, mdio_in, mdio_out, mdio_oen, mdio_clk,
s_axi_aclk, s_axi_awaddr, s_axi_awvalid, s_axi_awready, s_axi_wdata, s_axi_wvalid, s_axi_wready, s_axi_bresp, s_axi_bvalid, s_axi_bready, s_axi_araddr, s_axi_arvalid, s_axi_arready, s_axi_rdata, s_axi_rresp, s_axi_rvalid, s_axi_rready,
mac_cfg_vector, unicast_addr,pause_source_addr,
ptp_timer_format_i, tx_1588v2_cmd_i, tx_system_time_i, tx_timestamp_i, tx_timestamp_o, tx_tagid_o, tx_timestamp_valid_o, tx_1588v2_cfg_err_o, rx_phy_timer_i, rx_timestamp_o, rx_timestamp_valid_o);
parameter     P_HALF_DUPLEX 	    = 1'b0;		
parameter     P_HOST_EN 	        = 1'b0;		
parameter     P_ADD_FILT_EN 	    = 1'b1;     
parameter     P_ADD_FILT_LIST 	= 0;		
parameter     P_SPEED_10_100     = 1'b0;		
parameter     P_SPEED_1000 	    = 1'b0;		
parameter     P_TRI_SPEED 	    = 1'b1;		
parameter     CFG_1588V2         = 1'b0;   	
input         reset;
input         tx_mac_clk;
input         rx_mac_clk;
output        speed_1000;
output        speed_100;
output        speed_10;
input		 mac_has_sgmii;
input         tx_clk_en;
input  [7:0]  tx_data;
input         tx_data_en;
output        tx_rdy;
input         tx_stop;
output        tx_retransmit;
output        tx_collision;
input  [7:0]  tx_ifg_val;
output [28:0] tx_status_vector;
output        tx_status_vld;
input         rx_clk_en;
output [7:0]  rx_data;
output        rx_data_vld;
output        rx_correct_frame;
output        rx_error_frame;
output [26:0] rx_status_vector;
output        rx_status_vld;
input         pause_req;
input [15:0]  pause_val;
input [47:0]  pause_source_addr;
input [47:0]  unicast_addr;
input          s_axi_aclk;
input  [7 : 0] s_axi_awaddr;
input          s_axi_awvalid;
output         s_axi_awready;
input  [31: 0] s_axi_wdata;
input          s_axi_wvalid;
output         s_axi_wready;
output [1 : 0] s_axi_bresp;
output         s_axi_bvalid;
input          s_axi_bready;
input  [7 : 0] s_axi_araddr;
input          s_axi_arvalid;
output         s_axi_arready;
output [31: 0] s_axi_rdata;
output [1 : 0] s_axi_rresp;
output         s_axi_rvalid;
input          s_axi_rready;
input [84:0]  mac_cfg_vector;
input         gmii_tx_clken;
output [7:0]  gmii_txd;
output        gmii_tx_en;
output        gmii_tx_er;
input  [7:0]  gmii_rxd;
input         gmii_rx_vld;
input         gmii_rx_er;
input         gmii_col;
input         gmii_crs;
input         mdio_in;
output        mdio_out;
output        mdio_oen;
output        mdio_clk;
input         ptp_timer_format_i    ; 
input  [63:0] tx_1588v2_cmd_i       ;
input  [95:0] tx_system_time_i      ; 
input  [95:0] tx_timestamp_i        ; 
output [95:0] tx_timestamp_o        ;
output [15:0] tx_tagid_o            ;
output        tx_timestamp_valid_o  ;
output        tx_1588v2_cfg_err_o   ;
input  [95:0] rx_phy_timer_i        ;
output [95:0] rx_timestamp_o        ;
output        rx_timestamp_valid_o  ;


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Anlogic"
`pragma protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "CDS_RSA_KEY_VER_1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
iGDe174QOvlGg6aywFQXo7uWAhN4/9k0obvYWOWGusqCpX9dMpkOLvV7wn9pURJJ
SVc/k6ZrdDNN54sV3nhuoebBnew1pJT7xrjeSzcFzxk5klM/XPFpyB0LuSobaLEt
AH29AJGazQi9huI94TG7Uid9Arrcpb8c8zYWSAU51rNwORcwx6yzeWBNnYzBaEIW
3Pdv72fMiZwPyCaHLc6l4VLbXh7eqhvCUUDZ6vVDVPZdRmqR04y3M3R8e1LIzaqU
WT1w8/ICWtGI1T1T5KAUprM9gvKBqTlxa/shvKs5Iou0UTuWvWaWHONuz5HY/E/i
WjSC4J10hdZZX/ROXMGQ9g==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
l0h7NRg/On5Dx1GbkkoiNzM4bC+6eT9ViAio4lpYNxma0uN6wih4hhZ6FxApwRvD
/2z+8eIPycdOWy0UQi8jO7G1vIsxHrh/drjoKGuNW/afFzmuH6+W8erpvHj6o1vc
P6gVW6u0emiyfnga4TCrq4yZyriMaa8UdwM5pNVqnog=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
pz7npZw50nuSMdaeJCryzai6+SiicxpMF1Qh+kW4+9sOm2ud1QLskWgZuzOP3Zld
eDRuqoVvyHOrKEnNLe/UOn47reHUx9Yko7viXaJ3jVCCclgNCvPfR1XXCt9SX9pW
TCYnseV/NK2Hc9FTVJXaGNS1uzzpZu38P0xSq4q91NJ610RD/y544HU7C6MVDl2G
ZCMhdFsoCkzX9kbgj+iDM/UVbXpbDQNmBsYjF7MPr4c2LFDBfE4jIGcS+jPPOnbY
O/cTt3YySriwPCkHTrl/pbxcveVfetL15rgrUhbGnmCaiRIoykVRdxAr/DtrmB37
JaEHfnO18/zyeqy0WB9XVw==
`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
1uCh/WCyGsSf/cIm05faD9XOK4wtO53xOv7TPpCsbJehpJAk+BM2vlto80OkCl+g
30rCL4ZAUisOCxASlNIX1GApgHFDx2eA47XkjmaX6gxjAIw1OFxTfX1MLmEhqZ8a
plbMWGsLxzRQWtzXt6aj0cAlDiHsN0t+w4H/qDZnpCA=
`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
mVQwPFmqTyJ2Oii57G06nfEQmH03W2WbdlFr608tBLW3BrwGiZwaHyWMGX6kaUae
Kcc9fIH4x+HLZoFxEf65kWfFxrod45JDOd86Y/vNIq3anZ4smHca5j+E7DtqOfzu
mufzbJLWYC+i8+moWMoXRW9Lx7YtLkO/ne/dy5PEG4M=
`pragma protect key_keyowner = "Anlogic", key_keyname = "anlogic-rsa-009"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
m9qcOt5lHUz/F+lrpf6AiPTCWKXE3qqNfJG/HFNRiZ0nckVPx97nc4RMEMTbPAlf
9JGllIgoMFJ7ZH7Ezb7aOPNJkSQm4Bk5XljwMlN4C3xCMI0ALM9VstD55LiHiPF+
RlscFeoorMmSjhfzHHXPzK4LuaUOKjgOInTrRS6PuTI=
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 5536)
`pragma protect data_block
cUizKmd7oPh2xiQZDVcoDULaULo/ujZXYxisF4CZzEf3LAfghCSJUPUFDIpm1ysD
AwOpyOVdkwpsbHFBdKLyeHp3/ukdAcLGEZDnW36p50d6Y0AK/dBlEdov+EgG7/pe
BaZqenP5W6M3rNZFaTJNkPkPWBeul3WxihL7+bGa+uSpvZbYudAodr9o2dVbrO1h
y7FrhxuJD4J31Rg/vuDUGXGC/6tw23fBs7xlRLax4NU/eJTOBnQDGY/2jmV39j+w
vRbGlrspjQhFU7AGcQQDwLe5JP5oROtBQ7HjdikSfvJ+75Nm10huXCx6RK5k2wfs
qnBK0DvBRuj270m1kuOd+0PZmv6MCXK3TUT/Vde7PPyBsluigGCqOuTlBX9uHy3y
GBYSgmRCO9+QXhPr2tKcQDe90lSWI5igsXIcFPchS2YO3arEp5GLG9Lvmk35dIy1
O6pp7RrIIVnaxwkWtQw4gDsFhPOl+jX8gOY0f1mTimCIwGHFYpOXP+hngaJlE6w9
kO45jpKBDfn+9zrfJiuj7vpfeo8HaC/Xoivl5ZVGgpwfk1AdATQLkb4YkE7B3wZ1
nmJu6wmUFgMZUr6I1VqydWDOgQ6BbwmdvVIMMMy20EK6aCGZpW+WL/18aihYVaXE
8rR8H641mD01uqTqZOLvPNHuq30Qv8GLLRreRY/1grvSeZ9x8kE+07Yfk5IUP95M
vPnnSBwCj9U9P6AL/O4nDxFWi5W3sCfZ8Wa3XVvC0T22tiUOroZ1UyHvvP5NrSu1
4LF6g+6mvFI4TQUlazjG6PDw11nD6xjmSO17z3hsH6dkpEkwuMbMw1vJ5b3MbAjV
sxY8HCEnTfSEWKFrywMntFkdzE+UxZ80R751DPi1gEu+qdstbZdhb3SmjQn053N8
fsg/W+NVQMGYeOevxQTmztaw9kD2+SV+lILwQEZzi6Ks/TLXefC+N8k0vfumTEMx
3QC0wy+ZvZgSJOldaoF8qbxFSPmdOHOI02Rovj4eaRD8sbxoQh1gxe1egXxAzGvf
4OViKwRFn7wBUEBcga6f55+NHtBvsjvJQHJHxhm+pqEZm7ad8apvHbDdIspQwePe
kiROkXixeY6TAq796y4dhs9cpHJY3srE6KE71hPEbJ2SMtBqCifqFWq+ggy39qE/
TjARE/QiGLXhJbCQRDrAymMc98qh495L69Pg7Rqa1cJ6POVA8VWqMEZPUjjcCHJ/
4qMfgPwejd39bFeiLWsULxIRNlTEF1y0T/ZRtScX1aAqEOHjb5dRacUv8PRY0V0m
vvt94oAqtfO+m6AZdUm8FGeIJ97hG5HnEcUwYrm/sTC4cVNuO0xYjwvuUUZCLsVG
GVqn7MaTn1LTdJ5aETWzHBkvepxow5e97OC2miNducsLuX9KwJvMyTFdK7LbzFlI
opSpEBUxlLBVjTT7fTSaczZme/njbMcfFxjt3bh2mfYvejKeyTk137JJcvhiJtYB
otceZWaEur6/0lvLmtYjH6t2COiPMdpx2Yvqt04VRNNKCUdLDl2T+dU85+jXkJ2t
JPAPN03Fc21wl3mL7MrLSE7XD3CIJvgl3F3KKeWyc/qtavKL1ncsplXabz8pE7V2
y44Uq0b8ept+McuTnfelLO6DcPKpzG+b2GFMT10KQZ0frhPA14Lxh9deRbZA1PCX
pV8bAc9hza0EEwKu9JoR3R/Up68XbvdiO9XDtt2a2Ge7FGtpwdShL+vYiJKsIR/3
h43woopfyhXkggxnQL/5ChgsESy803Fc+ZkvAEXeVbKVDYUAdBZRr/6O+PyUFWv1
xqnZHNrRqfifTWiTkp09A8wFR9+vgWBYCqp9/c9hAURTQO8FxWLdrTkxCxO+7j+U
UhC/NgK5rfcCvwl3ZGiMT8U6FzOISspjbmXyUBdWCLD0an/yr1FEqY64WQJVbksm
oSXPPPCG/E0kl9jvxhaE7Ggq/siHBiLgQp+XdrBU64iuVq47Yz7H2K8PyIEb1pCG
5poK17cvmMuuBfftxeOWg+gMHORe63GGFus/iNUhzQzw50+VSzLPishpwe5yZsC5
4JIaMaD4Qrpl3Vz2fvm/7HxAdgvusfdevzf5zYJJnMJh19xxLO4FNlrEI1VRGNwU
K4Jx1AmS/QJKD6RwVky048lCQuWTbmA3uL0aHIo7vWinei/R0YO2oa7zylOMMArH
cZOyQy4QH5ee1UTV1UwTsBfA1u5N6XSZeFDDB90pPCmr0jcl5SxhL4waZLIvjQhW
aZrt4lW0J99CVQnEilQe9YvxKSwiCR5z1cQUWyH4o4NBHQMvG+zDTnx18mjeEEX9
8WEzq6FIvpOGe8j3hSPOvfrEFE8KMdaQXKBREWAiEVvqCCluDNqlqM3opCgAFt4h
7PWV2+RjUZgSQPUcgL1O4njMzzYC3zwzkL2CMXAuuHwNzl1JxTd/fmbXyjF9bZfF
c/4Xs4xlzHl7kPDnW3PEVkqu3CpcJ19SHYT8LqH/nHRUTdvz/h4fJV8pxZrwWSFB
vs8JGy6BVCK+BxzgCE1yuwLHCQAECdCxN1/hb7GmFLYUBR8HepC75Ix0CekeKXP6
e7L5zED1I6WQ+fy59+AjWTCBcXuCehSRy7HtrBQpVienRGU3+ECohrEIy868BhIa
1co/xV4a9BYxeK4eh7FZRzG5baz9JgZr7/d2Z8oe17wXf6Jg3eJ7W/yExOnnX0xb
OPiV+U5g1+HXT/rEJcpcbdkQ2BqRY9b7YJ8xE25rGIxBquGW1EQqa/gD00aAIHQb
zb9n/kkJN4LTmcDsDiiY8K2X3hZYCkrbMi+P3oCK4vgF6oOhuIJzZrG4zfBtcZ45
txBj43nPgsqxAhiu0YbElprFuRtabUitjhp827xLSLjczGTZMKR3EBLrs4g4IbVp
69wjTTIxpGgP6/NgVyRJrDvj4fftCeByQeLpt01OkR08HveuaKmWfz/GuQPSukmC
zJS6Iu40NxbX4fCkQwjBSv/LFLwsgpX2URJtnHrkLP4jpL03x9bSUehZVpd0iQO9
2dzmJQiqBDscCBuM/6tANl9TbiPxxTlWIPknFCT5GIx0wAyona08QNFW6dvQoD4S
nr+LLIOvnHqtuAzqELooEC9+kpPz8ta0Al/nciI+13qpbkzoRmdY5rqKnrVcpt0l
ce7NIEeW/c4ng4H/mUPC8tAdngvBXz+9+TshZoTek/Lkh9LVUUX46ZZsjK2KP46A
VaCWQ3YuKFWJ3Fe65ZLb2iTdWMeQfl6DOfEpH+RF4QitoiBLWNEmL8Oykg/m2aLi
0W6UICYnkHTcgHLWDRFp5byajL6ydq/T7jmOPhiQQz7m068uq8kO6nTN8NWENOIc
2iAcKk0j41Dh3ejN6KGbjUJKUtN0Ep0pC/sWT/mM1VXd/07EFO6tLHSu7gWnZtj4
zYStsuUBYVcB6Wrw2pOFqr6H7j3gTRkGX8uhCR+rPlQ45U9x2M7pWTYaREUYoHHx
4SaRVlVBJA8p2au6EZAbUIj3OIqIlD58FUWyOhxNbOW8W1q1F7+9b14gE8yBNGYp
J7U/5AgGuM+dfCG1Q9AOJM/D3Z9P5T1oXFccRIVL7Br/5iDeAUT8UtAJXs5KQWrT
zUd2+75yW5uyqDaWobH11t0k+9CxSa7p8hlRbpsQ2ro0BMgmBiT8qxhI6YOpQlmE
FpCOqTnRjiqQt9Bxw6HIi1dqtx7XHz6zxWrb/W6oRlUoYH7WLwQcdMosCWFvUG1o
y6UjsoKwS1D0+J8a19SVgb37o3eoeawvyirhZMKq41QXp8oyTCaMySSnzPP0cZyd
7W86C4YTAmEwhchaDllzBgAFgsOxoBOL73mBQezttvydMFcEJeHOlmWo5MYguCbx
GvpKl4ySW9ZzQilY3jpjGt03AFeQXglg/2+u0hkE7j6kzpcwoJqsM8BzhqwaS9if
y9Se/QHdSr0nY1vVbb3QjCy20lfIBWZuNANK58F/MY8rjGSjHJgm7VHMTz5Ea6Qa
rMuKB3EQOwtMQ+1qDEt29xxfD9fqzTWRJfxxZYgqYKkY4YmfGrz6oBcUgsK8Uq0X
UO+t5mV7YEYRlQ6Md4ms7kM18PXidxptL+eogRbJfWEMD714rb/C1scr0v/o9vwn
iX7hH0UMbf6pgk9TfCqL2pS5fEX8LZlLLjXjI+91BiITXflPJWICAx/GLnGZeeI/
AA01lBnI5pM9AhhfcU2bEmQsa2YofcoG0gaMNfJ/YKknTYGsZtptgJSRsrZiuUnZ
Cq0U2wZ/V3GwP1rms7pPZu//2YTU4HIOOYDZ6aLtE8j5qrLhfF94P8ve39wcnfEJ
nQZvHM8sdgK1FAx+t4gU8I1fG3mGDzdtjlkzyriGoaKys7tvV9E0dPBCN5XkjhtK
jxHQpS4pL25ZLtbOeIlL9QKY+E0WJmn3p2iBa8gKFiVT/KALlzzBUriLQ1IBEORR
K8goJW/I2EVQrOoi7UVlV2hiogvd6xMoGm/SWNm3u1XlzCnQubWsna0TUYFIG3YD
vVtDk0KAHqxaDCqcD0zSjJb6NvrDKWqtCBLCPULX3ee7HeiS4Rq9rp9box0tX+qM
jATT6XGagV0+uBiIWDALWCJTfvqV7bw8vCzrxehlw0XIyu3dyt9CJu1R7e454RG2
xOiDPnwa3WSgCeWVXEwPzIYWCD23azAxJmbBsiJfgTXSgbdV1t800jpPo+ZDjJ2Q
MQVdWdartcPPD7gjzCVZRoY+RjODjkEi6VnasE4UKJ8DkrlBu0ul+5WYOpJulRUw
rWnsPoMPTuIH8lLnvWRERHGvaHEXMV0rtg/QSbzlXMGWWoT/Detda++SBZCsjUeB
OTIEvfvfoNZNNQBiFR7rucdZ49A2XO/PKl2gyQbcNYbtVni2AdGQsGkvLQ5ksZw2
NqamXDeUTJ9qt2t/85q+UnDJq5SVWJq6CKztw+kZX38cfAP6g9hOynYy60LBgrVm
KfgA87Ot70LPDJ57uQWSFUl/DFR1/In6AEzuaeYDppvRwy7VUrggA2wYvM1g+ZTs
PD+G6hgRBSBQd7X6PSshBKtfu2aTW3eVgPCMN1NIFgIVtVv7k9UogQyxCG8B+D+V
LXdxjfyl04RHrSQvq9WDz5+/VtcIRwg7UU6r+BDhvIJkFTh7p+NjTGjabE5NFf8s
LKsq8It6aFiQhSQKH4SawWTOG945nBaaEU4jgZms8MP3nL6B5U5pGuvV9m9MAPJh
iCAN3h8y9W7R98xXqUYo5oSKBCg41CoQ6bhyWBr4Ml6VuogAp9Uy4jD/Etb7OGDh
6dX3nfJ85Qd/4Cu5rgdZwmmlWgtLTj84v3YrheaMlnpacaJnY1zZUdH47SLInj8u
kG4hqYQxDWuNhOdDg2B8q0lWkw3aI7tNBpH8BxiX/ExLbKIHzObbD5HOoVI0i8+h
/lS6c2uCtTYF4LRUuUba9vjuIOY9O+fYsPV83ntDwlyk1c+cfQ/Nl0X3xe5u5sj6
sgSUL+qf6SiN9cX4en9ajiCMDMK6H4h+Wxx4YHleP0ACXrFiY9DRqdJ6ePmUzGJp
/Y0NMB0auhdB6vl5GgYyKq8+T10HKJg4qeRoNtVUUJ7i/nRqjqQ7JDE5/UB3W+9/
txDiYlS6xfX9Epy8d/kjuOj7TaVUnSwzoG7O43cCLcoMSuU1mLfn/wbv1+9QLvaz
DTGm4Xx2TpgSU3DFRU1QBYg0SjrmscASY/q/VbogiOceIpJCw4422psI0wiMNhQp
VNoY01KtNYblruvwL/aVGReaimBxvZAMcV1SLA1+ABcDUQJ+z8Crpgw0izSaviR+
kciQ97F4jojguW7q7O2HQr65gVem8eoPN2/O4jo2GM51Xe7+u2+NPUu6IDZQUqdN
+eE3llOOY6UUKYNxzM3oMhn3vsj5+QE7vkE7z4FwCuC1dW+HGS18mkGgbjLv6kpT
LJZJoz8nMzkusNg4ZPiaTG2yTd4Yj8AIs48aOv5TnLHvqwyXT/20+NCZBQjQRl5p
Q1tp8Nzyygvlt7TVbf82gCt0jif9bstBWD78Ovu/2HjBkn2Q608uWW+XE4/QNBXF
9bxBOy1TndpcPKutrWiMs7ht3I+oVL/67MS2QcfPvq/CH8GRNQD6nlqyKoi8GNNb
2105ASpcXqDk3XEAB9C1KbrcrfcZHgDI8G9qT1jcyTKcKQq+kQn7nVupVlsu2mpa
8urMuT0Rf2WAn3Q19XnEuwCG6Mn3ocUMOBp4ChMDiPLJhgND6hqC6YoGYPxsWlYx
roWAU6Ur4mOOQaGskG6JFYUhVO+f0xsq5zJ1F5YuHhvVyOjJQJ12ohMZsfuInr1p
mkKFlFBwAMEu/kuJLFrOlTmU7OpY/V3/6vw3Ae599DZKCWYFFz2gCevZhmsR9Fkd
wJjVmz63vL2J3TFRcbcgBC4AV7bKNDZ72TR0G8pqYLWbVW1GfwpQEVxgjtlbNsVw
jsuTzi6dywWTKvmjraKOAj9WRlAhUbl66aoVIiT9LuStgDbZyhO88QxcsN/5lmYR
sm/dLbcImbOpCjOOjFHBCvb6QuXfMTsDZDMoY8tisYjokiKi1dW/FRlS/ormsSZ2
VVHN6FuHPC3yxSFbwsEuEhzLbVCy5mtrJfptZ1zt/dDU2R6SnYmX2ypRWagYYegK
pkOdfQQLjdJPtTZO+9O2hqzook1iBnQe3xgrOmK+KS/zQ65NWJ9/nL73fhOStYFz
WgTGSMVOPmlx9eCuqX7T+buZrb7aEeRDoYc+gmD6BCkiRJXf97GBh9L4tlTsb74P
/K94ecSvtXejQskqZw8hsGUDmPFZLOoBw+lQ0n2huU9GOQhEljANmLEOIJkwEq2F
X5WptLJdmfilUdI6GC8r3Xyz6hfIDfKht1zSOimKxaaeDHIkaET+15Jkz4Xl7+9E
TnVKK4e/rpHBnXoM+gL4G4IweLuOSUyb2piooSeH7/wLl9fQuSWjJ8rwFOhkUioY
HNTs4sRMwhHf6G5YYO11//vQkWdKaSFgcZaV7CVwdBN7NgdPErych2mg8Ay84Ley
tMWiYGkQuOGhHBlzp7YhZ4nHJFqbNpj2TEqjNJZSKyNouFVpcZp1gJ6SGIts1jMO
xSOYZe7cvkhARcGAXXIKvzHIctuiKjZlBQXetzoxAiL/G/w8OH2MYVPei+NV9jpM
quFw4xsmPkdITZO5Hfbkqyeujfv+bjT+4j7Rn4QRM7IsNEVhWd+jsknlqw4hw9Kh
Zp21W9vSsOGBpT9C5mMd0pdKtoO0C/Esj7d3Yak098bThKS+gqObzn0UmOYTfDMb
DSHFV1r938IW4rPAd9UgC3DB0S8Mt4jK1C4rueWio1FETuB8GrNhSm5gKMmY2Mfs
bjgWnHdvX6hYt2o9iCh1vPWsVpsfruGn20jvU3blU1CYOt4AwYkYXJCn7zYO14dK
462QxQHZoY/XmHjFgPESbA==
`pragma protect end_protected 
endmodule

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Anlogic"
`pragma protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "CDS_RSA_KEY_VER_1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
cbmGg1yiqOzlZTbVYXLPLT6/vDNIzKdVp+cAXtzKATDo1qqPwsZZwW0K08GnpHNT
kqMSXqNu+ko28KGe4/sz6sbJLpYb1A6KUDaUqNaPRdXjm7sM1Q2m5/bp+ofaSRuP
03CfrVX3boFCUrS1MO1nGE7YgIAuJ0aS5G/9looGyoDqhd3rv7ZSD7+sd9SQwj/V
RaJLHt9uMopUhuQSZXdEfyfZYrAIEZO2XOhN4XnqJxyF+nDEkRAGujDfuBijoPK9
ndy0ADQfU1qYjlUKaNypJm4GToUJPFmGyVC+w0x8cu6r384kBquCmQIzXjGkiBi/
D3298voH7toy5EheRhvEFQ==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
nW6+ihVzfoQpkFBxnXVeI3eCD3Zf6aPpmhrYGTMke41MAVrlnF7NGDBrYKpve7KS
joaaLg304yBlr09It1MVsa7x5hoR+uyXGuznPhvKsKs920QmYkw9XR31Q3l61IkG
ENFp43G+bt1/Lj+IkhdYaMsFaL9IYyVCZalxXxTFwUw=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
jMtncoOPZjlDBa3wOTne2zFc/eA404LlfePFlVdDanf/Z2v41z2uC8I6vkKXZyUE
sousX13rzpKZs95eVCpg0825NInD9jgSE/Qiai5AVd6EHqLSIUDKZIfiq5pIomHU
1T72YQWjG6+KPCeAueG1hDEKjoYADAQwcxwdolvg8FfrckdEGXB7XWCxq1MJskBt
MoDoG3N2Chxe8Pt9JXl7cBZ4m8WHoTjeGLyZOTbyJHdiymQmNCwPyN7jLYKpD9W5
CBsOkgU6jJK5hyn5J3QAo8qCje1v1nfbE9TsMTXI7jFmQ1zHfvytLEkdCUWTWFcS
HSqp8sHKKj30XMVrAv1feg==
`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
OhQd+7NF8cE4fURNw7fw2gP4AWDM+qQSoVhcOAnAdx1/QB7Pc+dqhQS2F94V/ti7
itnBXE+V4HrJrj/E6IHniVakgJylxk8gRjYR/ZexcOodwyvW4SKWgsD53ELjn4W6
YQXNAIuZWIZ1yD0nGC9rVu8uz1gAV0hd0L0zwvfG0wI=
`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
b9eIw/SMKFlbEJElLAm4haEyMwMVKrauek7KT1OLGSskrfKqUk5Gr6l42EnuTs96
eXyv0tW4fh4i7pUbsegsjfZCnq2KwLlrq86LTOS5QI87+JbvIDc+gwdSlKNZF7W3
2Vyc9rp9Mpnt1pVrqxHBtSHofNO783bfyM5WSquMRMM=
`pragma protect key_keyowner = "Anlogic", key_keyname = "anlogic-rsa-009"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
NxqCKW1wKktQG0pPnXpNk3F8TFS1rfXsqQS56eWnGTZboT3wwT0wSEuDA6meLi1K
TSh/bCGcehADrWZpf+hwpYL6EPwspsEywCAylg+neM4GzPZPrQCA0K2FB57ZVsTV
29FI2jbBr3ajpp+zSikXSfFDX5Sux3n9qdRNm4MsIdQ=
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 325280)
`pragma protect data_block
9wGI/m8Mx0B52Bsr/lOho1RivjyW6rcf41jLUn154A3UEI/IyVWhKe/Pt1t7phhr
2h+8qIB2pUSKKYoyAa8jJdQpDNS3Pwis/Fjwg+EuNZB7vPeEkDk264JUhx1GkAeM
E/c5M+fWmuDuUPI5F3PHLrew0wzwXm3mDWNtVT5y4pO5W5c6BK6Vmb8/8t4ZJRr6
RtTgwFfpbyN3DifvMWwAbZY340x5Nqsbpb7Wjy5WU7xcXxbpYdggxOKppNomq3Rj
DvAkQpHfThW0DSnU3G44jTvWPyWov4IorETUTV8Kg6DqbgxhBeT997xzbThTkGOW
/9lQ6mcyted5S9bKRAhL77qdolIwba0VgR65NN0z6P+mb80ABCwQ3D9Qe2/PN9U0
n8Uh5YT0v1HzFtcGD2pI+zO/e3v2gQ6EpUvJ+ZXLPfSyfPZUu9K8KQsM/AJqqIEY
KwYwJnsIx1Wssx18UTTllRlujoRsQAIJdyVXK++1HcW5je+MKoYyC7TeXTUwyhR8
yIzt9J+pfMPAPjYa5szoFNT+ZhFCEMw92fiuaa8ZYw/GsOsZBETLCUD3ziW6PiRp
oMxQQot9PEZFp2cPKFXvMfHMEZa/AvHtK3D3yD2raUYZc/Anc/DHyHGdABaXR3e3
Qk92Zub73zECALir8lXIKyUNud6ZAl23nTZNYgmYjktoauQ2bOYL+ZILAO2ipAnL
8WPR6PTjyqfOm9xZAm5arGyiISzyMuOpLScuS25ClBC9lVNwJNdgjfrYhHA4DHr1
L8RdmxPayIZjronFEDcBtwNUi1I/k8HE1k4b0PC9k/IQTbm411IxjBYbyEVRouR2
sUCGsbkiyUrONO5dVQn+cdrePx12EbGX9m16c5CQZ0hJh/WttoZu2yGmIOoBWL+I
Ussb1Ni7V5rMjBUlhBDIzRaX9qX/8n1FvFIMr6CFshbPKfZDwpUrMBgDJ2yRiM47
DvRcUThpiOKN/NNupa9AKq9wUSfXJ913AQ53q0SecZwwFyM9vie6LI1roCOiDNdE
hFNm40YavLCiboBbwZpXwS5dEKMlwLBcpgLBHzvMdSMs5HY4oXdJh/Ba+6nYd5YI
jo2XPZ8+WD3+ah5yX1fwXSWP9Y0aH+heyvHRYanFda6fw6NtvdjQV6aUTCDkJlH4
BS9kIZWpOhOEo4hEzQGjSjyvGyjEhUlBJ0FFKZczaP2VLtcAjkYv8DrT0Z3bk1iX
oy6bHcy1h2y6WjZ8Sr9OybZHReCPXF7NnmKxbkJ5KZS0Bwe5h5Hso9luudDT1khX
e4vTnjgvPvBD0W9bn2hbz+7wkPSb2QOPL01YyGGn1eTGxBFA7ksnmlzhaVo6rS1i
BanpO/SkqHCAf9kDeHXgslXAgWA4F090mZ8F2iUGOmPu1lWL2PLvXHwNYyKx/56x
QPiANwEfWOdGTC1ygh3hn8Nr5YLUP9dOCGXCSXkI5ywAZQOHQ4JsZw6FYryxAJQK
KibBKzfMZtRw10Xa8R3dhNXtT5v88T0boC7KJaRucpzzfrpqMuPkOAEwyETJUv/L
NqPNQe5aSulxsywGRM+d/qMMdXiJ1WChGrltZIcfS1jTY+qqO1XXDhX94ux4Ry4f
MtagRN0yFTjAtEvbhAxl+Tc1hbhKCqHKp7QTR9BcAbfiHP9f+pm76HxS16UWulPe
KFaJPLax2NcHNP+JqTohwjfdpgqZJNB6rXD9f6OOoeXBBnTnTgE/pTYPJFpMm458
3n5UA6QX9VwmdXzgH3zmcpRvkFSElYuNebznhUsqs00d868BnGSKTYQohVkDWNZJ
w8lwRK6JwwpDSXExlBlFEnDjTqyoyPf0HlTqilsLmVcR8l7v6YW6Vjv5Y6fH+yFU
ul89ly4mlvLMFhrivz0yLNvYEsC22vr95xzzHFc5skKCmeLPNa7dpxiruPhglmNS
LnlgqfR+SwBx+SprL8C1I5kzw5vlh3Ct9+mG+/bcDEjQmVUT+KNpozyLIGvkR1gr
/fDhBuaaCSjtLc1RD33ev/4lzgyukEPR85TzcH/RgdOL2PwcBu4b7XQJgN7MkRLN
iOCLjg8NP4RDo4qImN+659CsQHkZwRPkhEnzO8r6gZU7Rlc43T81kPlqFrrz6fEl
CbQX40KjhfgjTody1BHv43bPGuUewembe02mv0/gvqskgpwv6X+Qs/d4OBJRctgP
NWFAfjGrrc3zD5tJ3WByv3emqi0G2saDXm6TrV/tI2zkEYBKGGUfHe+cs1C5Lg1E
BjPYqz7tqKmMR/goVutwoW+rqLHNuI5/KtozTwI2kJecOdHPsuJpHEc8bP5H8n0i
yHJzmMeWCUx5CErKzxjn5jnh4tIXpUikANQR1ZlZvqcdOnOUROTssbFN5qrcMzqZ
VXAOlrD/qlJzGV0HwuonL4LUCaSSzSyoy2/SYE81S/iHw1DxDgZvDYy19Grjeu0a
XhiBunNXzupJKzaFl/PNsN+gY3ioTDw07AXeqSmN51s4x1k+DpFa5pp5jqq01PDY
rgB3rgWkY/GzcHnIHpnkQ8FuoZBfPyDozWA7isOwEp2G22kKW6Bw6/rUY+n0/c5x
zfLQ3gazOs2dfBNWLUxenKTlK9uQ4IPJ3EsA6W2/FBREEWz4FrzVY8UIvIE96N/C
XYW80+bCfGGJqOKNI1UqMsXkgT6QOLr78WkcLtahTQ3KDINdGLyKB2iE8RjcaE4M
Jpud6U1Y1avJlI/ig9VT7S6DdIfZOqj/rCOJmLCWXGZNrEDneIVVoQIIZy7X/5hY
TiNonU3Rm4IlPFFFg3uUamc7qj4JfVAwtXRfy3DdlecAIf+TRVQ20dGXJHGbMQm0
hHBbgOWhpVJ3IPJXxWHsrvtPlbvYRIBFXco7R8Dmv01faquJHUWL2yoBPMN760W0
yLDISYkuI4t2pxtp7suveLr24nVge6D2tgiABI+pilE+iEnjUiAWaE5xoyu7bnt0
SXS79YlQFXx34Z9sDQoeUUhyhJkvMBDdWJ4r6K7FMSpfg+uIfO4Z66MCnbLGU42V
bHlMg8CHaO5Q0G331B/kEos2DTpSzjOTx/A0H+0Ouv6P5suCdJhASsbFFroGMYXm
14UI5FT/J3tUXWV2F4t6EiwwMglUItOAdod36zM+DTsVTd/WSZLum4X/5QwSWwGP
Uxz3QQ6QeTsKflje41+k0rMZcEJgoPQy1rzIUEUA8UZ2UWOH5bhJjnvsjWcP7mwa
Q2PWvmWw1Vaa6m48wgVT2z5/U7xvLNO9HbZMByXP6E4RMcO5yudbTtyq9Rf32s4Q
5SX9bWBQtTdHeuh++jNgowRNzqvXgLPjeuMyiKvXGg65PZqOk5AmkUQ2aRoYpEfV
dPg750phBA5r6gpA3r0x3tRXhHATM9u7TJM062+Sw9654GPIHb/fGRvQ5lM5ETdf
0d5HjR7bSm8HcGVvOn9DsgW6zdaKrRUljt/a/jJOkQSxTn+sHsoRgQSDJ5yKhaQn
S/EVUadizCLbn59SrczOVNvYwW9cnPJfbMT+Kmq/b5a8JiZR/7OD3vsEj1tCkawQ
riagQdKFThVSxRdjGIKckXWw5Z/nTQPTq7Fbdo6e1WuJmzym8N6OQkEAHwkDm+lP
NBsTUMRaZ5peBfs1bG3oQEPr/k3Ga4qQwfKNeGYaHji0fm33c7nWQDkNSlu9T0DS
1dqnNkoHFwX98In/QkD0eKANGVQcC1qzl9MOn7RxcJtoyx8vQW5w8Hhnc3nFJ8Zv
uLq35F/w7Xg3vScESJ/8NXKCwUdpzh7nGPj8m4mPLHZT5H5+1ey/L0CAgUadom01
b8rqSB4A0HOVC/8y41UaZY1O5fMjfg8dCprH9VnFG3rBRMyYykQtl9JFWABJklA8
sfdiQ4CM3bp22phCDIFBbL+MddjKaztNzYIsvxlHaXJt9EkGm3RKXcbTuW5GmwBl
3l7MPkJX7whNEpunVv/H9UBoh/L44ZQIUwCn4zwJOC0AB3xVmFYoWcY1TPxMHJUo
H6ULG7Ui7jswm3fXwlPChSPCaeEKrci7lJFmHX/0rhU7U/MgrBYBYubpsT6F5HGV
SzUZswk0VNwULIui/jvWgkOO+hhlME384hDumjcqEno3UrcauKUtWroGSx9AtMpA
KP/LAC1lnlOU4As/KvGm9ZEpMCevQtXqPQ9xDQ117tEAFuI37/Vd5v6lX7zfDbRX
b4ZpU1KCEYPLbKbSU7c2H3MtqETpZ9dg5IpWRsKRU4R771i66vYSGcuCDAk2k+Wb
vxf5SWdJsdG1W9f212xxpdgEVFOpKhyY4YSLRGS/rKnaoIGcaKAL1uPOaLhAvrPv
+4BbxllIkJIGwRozcDN9Sd8lcn4h9LUnGkC2L21VVaEmHYOqqvAKFikb4oCWVrtm
yUDCn7Kso2gMhJ77USrgT2/WkIOpShABLKbJggrLNkQ6SzLI2UXYCiJmYo9hg/5j
4iIEkZOw+Up1FTry4xxcpw6v0jlSATuc1vnq5DLxykbCB2Py2NXY5btiTQmk4mrW
lagaFXsVU0rLuuymRLqP9AJpTNNDuQrqq6FEgNZ2grLyqoE1ncdYSif0PM+J33/o
asxHFVwaQ7kIGDXke5SvhQ88xjduNA2WEU5NegkPgnpHFQ7pHvB19o4exVd1lVy/
yShOPFjoZbfDwydNf4y+GQLKmC9LG1SYRCTzC0YGWYoNcuyYziXoE3G4FpJCdgo0
iOJvV+EjZ8JSUt/lqtZVsd8bdyc9wJVz+afOwarodevFmsIDbsucw3GBIN4YxK+Q
fPhZzEV8TuliAuJrbHvkO34PQ5iCdIkiSyf0zYOb9juM4zqx9nAxMOrGCjZQjmUx
DLp93jnvFG7zUxaP7o+ucb2R75m9KIuJuhtixUMLOlQwvArFFLuwQmrDC02Pjgjj
1nNgCR7y2wSMLMtI3WjfJDbaQ8D6eeMCwZ5fZ/7GePJ29P4rSOommXb3AuS4mZtL
HWDXzlqyl81pleIPbenrBeKlTMf8fqFlgvyQpDwO333p7b7mrVj/JfyIblHdLKZp
UfOVr2pmB7bctokXiaDobqidg3B8vCjCCzuqxbI5ClE2VVY8Z+DhJftfwZ66nZUa
U5ixVL3GiMtCzY2owX5z9LVBErUJKnWW0HHv6jlSBwazhnGF5DKuKy/JGa6MX0Ac
FP7Z38MtdBHbd1JBFMX/3/f0r0A2hRQWX00tBhYXW129Q3FxusOrBYit+eZlXpbZ
NsexbFtrabj4lPCnmcZ76RFcvvOYnDNF+fi4MlGoFifYOFeigGk6hMBcSEQwOViq
pQu9lNYrQZPA8hMW5xUKoWIWhwmYSqGtiWl9/aBjk5WeD4VAVICqQ/NH+lSHO7Md
94LfALjUTjSqDRgQd2MdW7ZA8O5ko+w/dwrHGaBZBViUwT8vfecqmVuYX+frms9A
Gbo7s4N+3YLLrCLM2ngL4U1ry2iDxq1hbLP3de73DeyeIyoUbljpdeqtZLgpWe4a
A6LSoIqkr464cJIw3ekdl0A2NFjHLw0XDg8PWMNxB9RHeOhPbChkk60AcMBOO2q0
tW0+ZWY32LxxSZkjxJgKnASlp+ihrvuH1743kuXWcV5KQ8YXhyndWPxgNCqpba+x
rhzWw8dT7ekW2QTmZG2BdquYgsiqH+XVdL16MAPJWEROSX3xzvTOa0Fucug2He+J
AlAQJ1pGZe6sYqwLRbeHVJOjwVzROSMU3nMTT59k9CTlEkZegvBwjlVGLdBMpZKu
gx816hwUaKjMmA4Ikchchkl+4kqQx+E4qlYO98ct0hQD2y0+wwMmCa6lhN/YIJBj
PrFRha3XGMFrS1yWUdYLe3QR7I/83NvGgAZscmSdpr7aiCP1KNZIRKpjxXNq8IA7
m+djIxdXr9eRZvkHhPEIfAt48VMa5h7oUgKZf9SXUp0RHMkoqxeoE0/Vnu6oiBVD
hXYM0+ZUbJAUQekQKZ7HsCxZY64zYL+cKOfiR+ekMZqNgghJ0RWXnllGuc8q+iqG
5ZD5pxY3NMuqeVX726x0+yPZq0d9YB0FefpW076dWeLuRXdh2oyRPIYcMfcxcWA6
2nm3qpRQfX0NI2LxgF23Du+GZH+rRgX3rxkWj4lLGXxcgM5eKLBbD4NoP1aLiWkL
IEGgIqJoZ4eXBCaEEu6cIhZH47UBDfq6ymCxHowJhofIKxghtrrQL+V2g/kh7hfU
BzLtNI0ROtFoKDrm98jtKsYna2saocdx3nA3NlPecUHPmacjq9OzV+FMsIlqNcA9
BK9XIGhwUDAKsIXR38O9w98htgwQyy8NpAR3GPtnKmrgBnJX2zM9AJDLR6U3d6vO
+PersTDR5qesVQcQwlsfn/4gZWfRINp/iSNi+D2ZI2g8sOifZogNbAOBAZIaJ/PA
MYkDSgXTPIb6rsJWf1iMSJCP/WpcyZYGhDnqyKmAFEc8eDVWUDUBHqEXKa6AsNqk
NmzKIs5XkmpUcWwqRciC8Z+lheSw+jFyzCmsU+qMOOmCgcTzPID7LMh1oUR9kAM3
/D3mFPamKINlbc9FXJYEZNxRS5ENQt6YCEdzmscxB0Y8eJN/50kbOhsLrCo1tqTp
Q1CONBhIkizgXUnFejB+zV1mJQ0WK1OIq3qaDREeQ4VCIk73+FU6IZp16ZRf14KA
jVXv3gWjMJoFRnzeMvP1Q7XjdSZGI0YVCpEE1WZtUeBbwAIGYEoloMSs/IYuFuk0
SZlD47b0CFFvpsmMq4eCQ3RqmqVbNSrLkqwnLQJwhRRiJEYCJFNMJerpg/Kso65n
c+kS2uh6+6PB4ufKtcm25D9xIVZ8gjFSg+eX5F72Yh0MVdCZZ18RojxH7nLqx9/j
8Jv3A39RkT3XJqFPNgYErxIPtlMm3IYKOfqja8WyC7Iv0TFZbE3rsNzW8Bf+JRHM
eY5tt2283ZYk4LVy4VwVdDm0MvxQvWLaKBJPRBOYscv//eiVsyHOpgW0X088hTEi
G1DfLMkLlRSRnL/UcSX5n4WWJfMm0z/XRwhzFU64WTUNeY2FWmxMiW4E/tnAqCkv
+QnXV28TWexllaTBlN6YjdYDios9aWWcOP012fAGq/qb2qhV2gZ3gVPpTi36CAw6
1B5mPaNzzplLPo/9U9UprroDq47Y8UJJ1lzs63r4WACKlhxDQ2lF264qVOUo/q7p
F9GbckzMFyXW4tkzoS+9H80Lcg5mEp5vaGw/cAWxB0Ef3NemZ49BA5ZxRAG+Lmnr
Dtqi6PVhKt3M2u9WHQhESUEYsd2dr0Hp6GjuLiQE8+vThZfVBDDYQzuJnifkqX7k
n1IGCKF7k/XNalO+SC6Vl1ARsMxa/PcpDML0Rk0p0tw1Jt0df2zilC+IlZMUqNcY
kPCHVsNFFuP/z8b10Z8Cips39YmdBp5wGsgPhtVE51XmyCoFLnhS0Xp5XIrQ8+BP
HnEVEZKgAZzXch/v/hBAhD612dEV768lxs8G4XxiclmGtUHhhVL9Jxm8oBUtB+PX
CJoeBIvpV/d5WddzJ85srdYzN57+pWasgXuBzxcivd4ak4CJji90/NfS5VImxcqn
5VTTm5clZDj3UG3btFvMdcuRcwPtOtef3wgXwIs3frvthNagxqkiXx78gKmoPpw5
x8H5Z7BAaFRvCQk3yPM+2V7uvbGy1Nol7p7qxw1zIoSzWq00VA/FrbGOzrqbEChC
1NFfCSn9+eROlgU9c7TQKT/4ioPX/cCGQ+En/GTEF2vQnEcMtFHg0sENa8h8g87F
rrvWk5SSKq6gXn3WihOm0rgAlKLGb0oDz4eNAqKAGuVsW7N7caBm0IzUSspGZ7Px
+iLukQEGF8Np4OQ7dCPfAqbwKEjqWJ/JsKi3BzHFcK7jm9S+S70LkLzOH7NVd23v
2uEMId5ygaIWS8ybEcBoT+JDY0fv6YJllbgKjRq6fsWhdpY1ueXWN1NFbGCBvP60
QjxXm6nt+Dl+MAKHVSR+O/8hFQF4G0WVlgskQVgdo+RAcnvnkfOPMnynVFNhu2/W
3I7f/y4Hu1Mn7tbFPYZSTja3dwJLmsuI1W966yxBe5hYwSFHDAC5DWLAKKEfcLOB
6j/IlLsFZVhCm7AhESGxn4vwQ6W1SVXbBn91/Tw+lqsDhUDsHVIcFHt2sClPmKH9
rdJZf/Q0PSuJVeWaj82HZXQTtNf9kzlf08SiJ0CnhUhvtCVnFZuhEh+l0uK+9laI
fDKjTaRRTekcd40vp6L3bhWX4gcPlKgGKcEdIM3VEmF1+ZAysV9zuA3OO7GYJPm1
ZDuqT8c2nvXq5QdgonJRw+HtnglcJA3OM2FoDP2cKDYcujYvYGW+8XLI4XnuaEih
eiHhSLW7abrHtR+TvVVC7/OOUlPRLQ4inKUkt2euDqd60H7tVRh/a565WPQmdscs
TVd/miovf41u4HCtGf5c1xl7+pH01Xdcl3wl7yPSlPjAmv5uA+Clxa2YqkpvFRKa
De2VlzrWfKx+WIs8hYOw5X/ooXgNhotD5wB6GiEkgoqM5tsqmrZ3e5diM/C0S6Of
LltY8+WdlHBnzvAYeG3fki9tX0hL1jRgeN0wOU8KXw5/c5wgznJLnYCMJiJm/6E2
txYTy4/FAeqEs3fIoPYQJHNwG0Pe2+AeWODl4aqGb9vTwcpmWUiXD+P4szV+fDhZ
0zOfMJ7LfdQSAXlWvA8KV/4MN0qeBo8uLXJQDcq6DZHxGvU6cQBP/GSbKPqVtZts
yEuSuT9HQrBU+twZdv/iKC9OCxAWl3f9CXF1jp7S3ZwqHMTyn/RzB+pbQARKBUe3
EQ+LWPHCpMp/oPXXxZf2Q4xDEBkDZQDnf8yeH2KwLnkM21JKvlytCN7IAULuuDDu
JOnE/Q8zGqWt3HchR8z3qqqMWr7gMSZldom3ZHfUptdMU5vzKkg9FacaOfJC9bZD
Mv8FPDYjR9WpDHRW5cCe5Ae/c9IbYaVKM5F/BNllqrwWHcBmwjNWkvd8iaxmcMCj
ZbvinaCuAQGS19k7XAq+b0AmLtYoBDIPNRj92T647CsXtrGF0IpIarYbD2h+mDk0
c8HteUpqtAjM49tqFz6CuWrTTeOuwqabi1xCDY616XX/RBYp+ewmZi7q1V4qv8m/
vEJ5HljxHIdQ6h+RcPmrUIeM4ZMx21JA2slCKTFvLfgYdKDNtBbjjEUccRi2ZLfL
axDXO8P92jcFSZrU0X74Dskm75MqlYmg9X/wdfI5gjvlQqSdXqVx6xsVsEdXghcA
1NVWvAS5ktiZvoHpDxw6MZHw11tB0sqXPxoE6ckYJLPEbLICk8zYwkdlvUIiYuFa
ep2HliWPkP24XqL7QXC9H9WDCp1rF/d+8ra+ii+VPq61vO22WSGXmTVhcksq8yqH
rxxDyBQ9Hn705QgZPk7n0nePbeG/hXygopBWcpinLj8l/YhvuJYe80LoCGyCTPE4
aHs0S8VMX82tPtHG2gb0qm24nKY2OixcqR3LvNxfp2lIiOxuthWUtrbuuBv2ZJUS
kNIBxne8JLX6hLjdc0EFSXDNJrbi+KZ1hjWXIkX2H2/9CY15icxCZ20I3y2U+x+A
tDOuZZilUumlBinGAz+2yIintJ59Kw2poZ0p/95DJDu6UgDV3D+p8LatpVtUg85W
WXNRExktjhlIoMTtreXgL6wn7+1xR3p5049np47H93jq8c9MLRDiX/0cTBP8SKjd
o5NDMHN+VICWgOnPAlDtkyAnovNb/2V9TGFdsfxAgSoODOVqS8Qmx89RtORWm1lP
NZvMZfeAnTiqEhP9BBm/eTA+UmzDGuKD8M71Qeno+uQNPTgH5Oup0T2j+RUyIon6
in5FE9+2k8X9sljsGO5nWZuNm0/hWCYE79sSd+2dAqMDICPreQm9NojSlGaR7OH4
Scgqi04WNM6K5K+a1oSWqAxMgqoukdL4omaR+pDO/qPExuOteX4t46HQSg5dwcVX
02mwELa5ddvcPHvA25QY0gpBGKeQLJgHVi8C7KXLN1FSvAguEhk8Q5lCR9RrEJLb
tMz5YjQkyccivncYLVoySJFPf08/beLKTvKAmE5JNi6rwMvDb0jofrpO0IO/Y+se
Xnlj/57wCXuS3Fp6Swz9ZaX3dJRn47PlQ5JwX53e4EDH8yBQ8exbaRp/sq4XP3Zx
4fvuescJ0TvNV8zuErujl9wWMdIjNOrEA3qLEBMZni+z1V/Q5IQBiN3oPfuJGmjR
E9uTKaAqIJBPnANIgRAxlXLAxlnKB3whJ3h58PHVxqaPsXxTOLeHk7ebsoXFO3hY
qhI7mdRP/A9G3XK276Wz1ssjnqFp0ZwWEnCx8+zdL6QiISbWj3DtnKz4N72aaapo
wznDe4xnpALYBfbJD5Ym+yBPcfIzzQEuWSL5qv0DxcK0ewe011xiIVpmE8VbGCXT
17o49d/UETzS3hFImFh+/dyWuvsTrAJX7WkkPa7q75z0C3GUQONXi/FA6E93jCa8
LxptWvirB+oP9sOz4R+avcTtwdsWOfOYvizkmvTGDqXKJVr4Sp9+BJyecWvC85oS
B4aYH7d3O5343xxeuyuMpF4zDa62P5tS+kaSyuGnylUMEwofHsBr/JapHXUW9iK+
1wibNRo0qpuRdQ5lLxMkSsXmLw4y7o6iOW6itzkyZQAbSSmErYmpc0755J2ibXn7
sO3WyRtWRI+ovnWOyBURyv7+86zexotbIINVpHPNuwdqX0DRLLf83g4hiVFSUHwm
pMEkQkW4niANbbVWkTK1JzP99/r7kkfADMhU2CQQsY3DJ07ScF9E/uMLhxOJQ1i8
qxZGUB9pLw97aAt8001tFpNV1D8BpGfhcYOl4l9krNHXzca6dNus82/MNqJCJFR1
Eb63RmsQc7qylqlGoi1Zxu0tpARzzDCrHTFSfsSdO3UjTNAuhR/M321U3P8a2Qvr
xXwgocl3NNw7jGkzluUEf8zpGqENWNFzRN6hsm+uyvfVN1cTFCsCfNIgBOpZytFP
h8ed0p9kxC1YXyjf4UYX+2xTDvIkBotwG8HwYtM/hEGZf4MCAhOnBkPKSObSTJB/
sLDIHEQE+kg+LQf8NnoEqA4V0N5y0KF6tLo9QSXXBvURZ6Q0prp5wJzmvQJ+RiYu
Di/uKtynEgl7tm8oI2XRxP9LPlJjiRQx37Xfta5aSqcxDZcBXs3BlFJUpnLLNhy1
sI0CMAXz04pV0TQ7txILH4Wg7irBL+jVyRqIY1/u+qNIGNkqDMfiBNOlETnHpIXB
VpzbaloiQCqXnUUUmkaAC96lk1uc2rHMMDG1OqdhbCQbGVgUIVTCeW1TI75LgYNo
sowvwmkKJxRaGix8Zm46+h3SQmpthDMMrqVfdm9L+Jrc8n4nTNoLRW4GluIFI5Mc
aMqJuQbdbZYkAybKhvRpaSGjf/XCStj+DBEi1AYcpuwwa/rPebXvSULaqFbl5GfH
FpWLBlJvFbRxwgMpUC1o5awUESVsuaSfEgguKVduai/KKv7AmmTjaRRLRCvZ6IqY
tksjDco/f4ZbNFQEaX/LN/9d/Gw+bima3ZTGpIc1Oseg856p/YDXbjEGHQUInHjO
d+sB5EdCfE7C6yDETD+KaujYvdAztQuxDFajojqoqL3JVxD1D8NxKH6DkTLvSf8l
9QBxVKlv2dymOB7hpr5/iwcbD0iIglF59vOuvzdAH3YQcLhI4Z0LjpxA56IJR1wI
WQKJlwAH8Z9PbKNdmqYzoyjRxGCusTKryDgZXlrvR4eTC5Dy3SEiIwkmLlsqOq0d
oqT1c63wBxYXYp5HCpkcgM1GYsf+BABiEZyh/ovV/iFWgnj/2oxcwcQgj4/vO155
KSgT8/Bd9/09U1nTgZrmUqLppJ3l50klQWd00DH2HQvhPMiFPBYlKelvigiZGzbs
M3mLWRnFffByrPrwtztcZCqsxC7EsoXiEzIuWdQE0RzuOS7vHrXFOLhNAI0DQoKE
LDt3w5bEt1/G0vr//p7J4JdSgPCitIdsHEwlCuPv07vY5VE42oEZDAzhxVpc0qGe
KQjIHt0S6h+9E87A1LB1Ok1Xr3eraAwB/ltJSCyUQqxByECe3Neezn3hl83KLQRi
fEY62MR9nX1QeaNygswtKS6WXzWOdP+EPnAIGzGoJP6tlAFFUdSqlJa5zfvZ+krm
hq+aIKk19oHr1eKO6PauTCJimrwSoCId7/1lV1N/eC22vwlN34ryyV2Bo4Y61mzC
G2gNRuRqVT3vu5hIolxo9Plf2Fa1EqjDFVCkZRVm5ke144bmU+xYB8GkPl0+7VlD
6NAVW/XXTgkqtWK8UFukeBeZQrEHwxzdJJnUU0FeETbLS+NBSwWqH0yY3KEeaEhk
ZwZ/JqZHWiikAJgRioCFUQgdFOG+cqB5oAp+TzMRRoQC7G4MxYLrgQ8sKwLHCVm6
2B9hTLjyy10fE9tPs6oZwlRujzTSQNKG81JEZaEGZ81Vl+V0i6U3oHhYXvMhZV6i
PQq4aO6BqQ+kVRqsqHyxfZ+Guzjx49fpm1EFXRB6yU+Nv7lnGPEw7l5RWi3OztFf
9ue5AXGhiZhXqeY8r++tOj1V2yUyOqRvndbmC/c2JKQWN2wzmqkWp3pCgDO60OCt
LZwn8prAzNLwHmK8M2upULBbOIe8AVafYkAvNLljsh+af/RAFzIv3unlXE78BynW
wjA3AvyhVjLx89Pwtt2l3fnh0d4DZHrAz91fhaiQAcQ4kauFymKM2LuTmxO+65GI
nNLpBNdETOZnQKudjdufgCrCD2/4QdLLu+9eQd0N1W7ey5eZwAPuJlEJ1LjYOmnN
LtaLm/TBvVwHkZ4Pp71AC25csL84u4Jknm9vPdSwxVS5VHdETKtH8pTavKNXg/f5
PwzjJOt8TS7zGtt2wr+XDMCUzrjY5oxnm2KzjzWjgWNysgPa7fIsNFILYmtQFnSr
4bRTVoV7+YvUeCEkoTqZxfERfi9x4+JJx8j6K6Jmo9olHKqlFNhmrZEEIcNrHICf
qThYFopP/2ftxdDpRvqABakaJ6t8ReuC6a6D5D1UMlLJAV+DjsJ/EYUDSVTExynT
iCut3/1AzcKGyUoJl4Jyv37/ILb6OBb65swNa830SesLdj/GfPh/GhaVxABpoLLc
2U1xS2xCfiPIGpgyIA9Fg/gN4T+ZikBztEyVm+DebQWfXydGTB+K+59tgMZMIXRA
yezObyH9vKGLFPwohQYhIwQ7mmLr3GS/zcnHy86aVriNo/j57/vwhBW5NR1A1xna
uRXbiXZAHnMODEL9JwpV64k/64Y/vVviCYCB4Y5w1Q/eCVa2BA2+O2njgw6Z4t1m
ALp/ne+LrXb3bCLy8uuraYAs3OkwI48Kz6YF6gAa99D1q2F8Za8C/vT7CRV4HEwS
GmtEt+OCFvUC3+c1/R1Cv5GCgNX2sQdmalcNUSEk4ETg2fTFBZDml98jYLjOuiEO
inG3wesq62I1TxBMkK+rJ438GWVyMio37xRw1cT8aOQhcmw0rWWXZ8LYTXvNfhDW
YrWB6bXrpYADPYVX7Q5LJdcobDW31j2HObuyzwHWqcIM0c6zcuDY7lcOccKp71A2
gFwYJkoCBOpsbIRHv0dJ45KCA89fepdf7vs0SRnFT8WXbXJepo9Ert0jANrJl+IS
UkSc8wKojbjGk/x4hfpUrHmow9Z5gyGOYlzPcm1rYMC41GNlpG2j17KdPHC0z10P
QiwTxdD0qDC00KNVVV1RdBi7P4pZ9Wqh9gH1g4HoF26yl8MTXtjPVHGkg3/SeRyF
w3Xax7ESGDYZ97j5EC/PTsgTs31UtjpMA9bRgxQi7gutQ1x2y1yCrHm4A9YoJicU
Eaf2c2PTQta0McrIMaozDx0Xpleinuq1PFdTSqRrP+Lxztbek+pvkNu8vVRwcaX/
ZnutjocUgJyPZk5a9r+Fpaz27ZA4MPucri9iET7M2SiXxSvC6riGvWNeeyOhgrm2
Hkd4OunFplR0E2BBjQgB8hLdps06ZmDO/YERCcEUXVbdorucz91tWYJAAshHZuHT
ix9ypNgy2hb4UM+RmuuOAYol0wUeRq5souUI3AcwYkLG2k7/NBDC4yNGlsCmE4uL
Kaq4q0aB461Wo2VBb9Tn4eSvsvMQ/6kTkacmho3hHJNYST0WtHk/BvGHkOE1VWw6
RBXrJECUxy+f8TId7hk2PEuO6Op7AW8FHcLaWx+3QC7eAdeup0G5MpXtv9E/Zszu
B6hP4JKuLC1AeMSbeXakEORto4htVsjfz/SgkGnSY6G4Y/r0WfirHYdKox36JgeQ
lD/b1pOaI4Z7xsXtBy40ynt8/gAZlMJWVxfzLm12IGWc9hKYcKWcdNvQY3YTxSjH
o7B+9d/w7YiMb/GoCSjEmtONwI0UgEhlPBQJ4E1pIqFnp8dmjYz7gyoN+7c5Ee7q
fQsOmd78ljhJMzEQpri93lNae/8zqoNAhnXYXiCbzyVRM5tJZEwzVeUNFe+HYiym
OO1O8YccBHOyjnLh86u0XpJiqW0oP+iEOXACOkCCHZpFhaiATJrq/+lTtspCEU4r
YPZDdPnlNtnFYqYhCm3zP/ZW+7hJYeBFOyyTPya08mnkr/i4aE5xr5uOhrjegknS
jDJab/VmfjBcUDAkvTYO6s/+ZAlGHJ+GYt4u6ZCrATqz9twjD+vha1dZ7mU0XRUF
3WLrFIEJvfdB/fKVxTc1+BIQb3kea5foaiRzECbb1RN3SvpCxrzUsuG+A/ysZL+e
wlDHWcEYRQ0nl8miqUaDar4YDzPUGuc3rb1o3tNzNoSek9hnToRgtcH1UUb5uZPj
GdwwFzegGjuhd+z0WGqUJfZUgOy4lYSEcx52GSz2vZOS98VOiQrdUPtGB8PnqS/1
AiQ6QhuSWtatEDVSyj1cwny28RhAN+7BACNlPWmsUBz1hylNO/2MGJr7ZiOFbso1
nWA/QXDFdhe+JXnW+kiKhZIx8YpteaGZ26UIXoIlm+bETDtEahcJ/rjpKbHbbfd9
XHhwpElqOG1q7Xba9P7/Jcyx+OqHIRRCjbdQ+YXd0zxceJLHXVQsRq/4c2WZVFZJ
tSwnkkXrMXe4Fvsx5FIUS+d2ymTegBqAUTlqc2i7YFxWUqk7FWuAStz3xZG3iJFy
jJe7MeiWu08cTO6dZ69l4lxXwwX6dQZKB1XODvlCL2NYr6v68bKwK/+l8Ca1TIsB
iCiUrMiGqbMZc+fXniMDsbCKGPffTorEUIRQ/3pNmaNejVsr5uZjm3Zi2p7vzO4V
EDh68oGzZoJio3DuqSYi7kXxdfn+jY9FwY274XXDddflyV1yXzeuN9eytEeJP4+F
YtaMuGHfdWeHsc5IPHGY9w0wbW/ZIBYEXrZdKiaT5/BXwLa/3ElYw1nHuIo5hA/A
5n5qV6uYNBeZUARjok7+Ak1OVktONJLqqhrqjzQT998fpoKaY70DhayTVJ8zCr17
PthSUXb8oGCy5BFc1yl5kcE70zRDkaxFwuCXTgzNJS1GsgJ94pGQFXOtZ70HUt6M
zmkBRbUAO7HnVLS0VWVyXDKHHJb4XPxKdKSWW4vi1xNmg46QhJYXa3detTZbA/0b
5dAVPTX86Rzbtyey2jGS0zefI2SLKyuIR0IU0h30st5Y9NBUWaI3w+5nBISfgNfX
CHls1FqlHZgaazmGto3NhIi5OMmYv9uEx3gbHILKdViNV3s2Myssadb6+O8b3cJR
8uAVlBUpqcIN7AkXHSz6s1VGqgNEx9XUtv191+wLj3u6tlwLtgLP68HZSxAAGReI
ykCmkxcW1wc0uBWI+E5iWMnWj54+VtufONDamm3TvVYizMUZcr2f+hzweu9sQFxE
KWBsxUzbTdXZqIMR8fVMBLTXK5+OhRF4QWN7PUK2kHngCdNBpx8p1NlQde617Bhm
IYO+1jA5OhNfKjRJMewQRXSSE7PKKmQoIUPgv/ZuNQHjNNMQOdZFKXNxYER6uA1g
VFvY4rD0vUMbXokjHXbR2ng4EhFTj6ceBXrh/v0EYsvS7giOxFBpg2mvY0IR/eYd
gtxQKVBty5bqQxug4bo1gd++cGIyVeQxppVlHEPdPclvfkiUL384sQFjhL9E+13L
muiMdNigqKOKNwEB+MfJvJGcEtzRChAsWldLUbGpjzHKz1OrJ8GVFdaZyzLoVDrt
N7k3pr0dpHKs4gKq8ZYj0qtVc37Y/RUsYshHpC82L70C62msuUWTGUEupDDyYnAA
J/xaXW1+6UNQ7yZIHpr6tsLtU8Tan4yXAvGCWhWabZy9/CTaBw7c5k7YPnAnT0SZ
IIZhE4weP1PNk7Uw0YnOS8uqO/6FH2Dk1SDwvRjzDTjynP3kqvoSSQKfuulBs3Py
QafJnfsjau7TteuE+1CZhz7jJxMHcmB7yBgKtnN+RG3E4PvuSrjVZctqr67Xuyna
fSmRbh1vGJC+4DtaEYNIFDS+f7f7uclI+y+Y8XX1Npk5fZDCpRDUR3wV4XVed2jn
Py36RMmHqpDP6/rStt8Ef+7buW4pHXu0+RZpG3k+LHtQX9nFSklAKxKqNCglHjpX
BXVfj7foqWj+jR+mGUXYsRoJDcj6j6Kd4toiS6wtGu6Yk5oMA5yk5Ne8zIbVgrKB
OPNZCNfJfdq9+zA8vMHwyDrBT67xVyukeyi2+zUhLKZcc05H88ZdaTnr9Jpe3QKN
84kBBbcEOQJlSCeA1P0Pad57gLYBgZTk2d0ljaKl3wHQTZ+Fr8L1PrDOcngLoChQ
OgGJBr/NrtZYVFJ040U/97XE2crqy/Drapjsnxc5oXWVCRdxz19sRRWzclBuz2l/
qH5ller+lQwIYz9qHnPxRfzqPgmUl0daWIolSUlcjidrZfXao++oKbumz0RUUtXf
HAHXNZcLj3AwyUmCcTBH+L6ddPlarSLfUVUGzzdwDDKh8+O1homCCzvfMfpDvzYZ
rVpMM+wDLl/5X6jOLb2YgwkJtf3uNjJdKEHMW5avq6KzMOLCd7XOrkgfTo+OeE4L
tEGLkxoknmqzPFppVLt9Wpv8bxX+nDUETnGzFFKRMxd8YHh+94/Ftxti1O9H95lE
1KOFZen4Um4HeIvrqjiEiCVtRYkKsJmU4MpIGQdOOTLlFg3po4f1iRCM5be0ITra
YudWw3JYoU3RHanv2dKo0VeUx1+moA4j4Kcj42rlr5Ngag6hz05TM8TzAQctkFx3
55AlBCLY4j+aCtWNk/vcNM6FeWtY38FrUU6hPw0VsaLn/m9hyrRS9Uf9DF5sCP+q
PEiYP4X3zg2FHPcovovasNqkx9LuBeFdUQIeS72ITUKE3fKkR/HTbb4XmCbcwSB0
92iPhrJOD8wyN71Ksr9c+LQ27uLjNQfSzjydoDdESwmz0hx5Hey+vvezFSYuSCWs
l7kceJV2RJeCQtrnkZPm8/DLwwfe14yly7SQCpZT6BVR/DVZXbwWX7g8q2m9lb+v
5thaUsmoSYEJdj1eEc2PoqqaUxWOhuIs+2yYz8qjRqVQw49xW0y8F9vdv3hMLZpC
G0e7AR/XW8boHKKGg5zjdheurLB+GWdaI9ZU8wm02MvcaJUIo6LT6Jgn82OhbiAM
R6tBfDphHJUE5wcTWXOcID8YRtWI+EV7vkR7VpaQm58Hv0zJKbQxblX/yQYIlCIb
iZ+w9QVr3nrHUJyxUJbiNDfIYEv7R1iZKG9Rew1+W3bI4RX06mgVRrkhurrQbw3w
4QkoF/GNZQ4857EmKJjUlEwxbwcoHN/jB+3fyj4mB7DMVs8wMWW/AktgniNAc+RC
tPBJn1rbmsukwexn/Cyd6gAJHCSF7NG/uQJyntoWpMOUjsm7K4NXyIOAQy577GwY
Mk1fmt8sSSWSQ/ezEh1tewNMx6wqiAQ9ds9ubxq9tTphFwpv+5zyIzk4cY0rdKwu
tMS5OuWbWLPl6y6ysiYDUztiaXi1tXBUIaOhJBU/kfv8DcUvVt2nxA/TBHDt3ySA
0dxmbxo67vEPB8QBR1lyVzZuaxq7juEWCB7pTQbCttAjqH0SfkteZYQuXvkIbUHX
zzcTh9qsMwj28btrVmSNSkthUlrmBHup26LeoKuIgxkDJjQAfvKLiH4jVrN8ic6v
DXuSAj1rG0ocRQvrbReLYPH+NHVXoQ4YUx8pVxmdfySZ7jFuUGnZ+QdKdgAln/W9
hEH0y2ntIw4jovEic9chSu3/O3SoIA85qKwhJs5Ax7V8OAfnD7F2P8GoT5D+m7Ev
bF8gRg1oAix8l3jBScVps32OlNY+24RVUqqv2giG6vGdZFOUBzJWSTwjjR+cxZ+N
sKd7xejJ5ApRPupeYE/QRDr0190BeaGhiVX1Qj+2NLcVW0CogPnmcmx67WJlBDIi
/woMqNrJG6Lg0diei+xGI05OtULwBNby0KfDtr/qdmbmhHi+BALav/2gikR6LSIo
YNUxjnzub6JsyQ6rQQq/8O6YP2EQsCnHmAFUstoNKk6PFQR8ICZNjMyvkO/YbdOv
UKTSuKq/YRWQPrgeKGt9+D4nIfi3KIIoiP6POL4yvlb/kudkhV+2QwLsr+REjHcL
uXKgrKe5GzhCgbILjzWPQKVLDt4g5wX1wgkEiSZo69wRqvhsPHisOm5A+9nlmIvx
ryT02K9OneFXxUtFRXaUMDhFm5GlKgkqN4k2g93FsVpWYSqMTf6edbtoUlvoN4CL
Y3h4WmC1O/gHzy9+r65TT9Pw5jw3Rvc90/NCbGbr6zo/wn+lmM9i06ySf+cAdwU3
JXrP3fuzqBifYdFSz7PNzRZJUGYFWVZBEzSX7bBfHGomoc4QqyCXK2U4M3HVTbP0
JMmWNtkk8DwlTwJrIv9Q17/KmTlCHcUrptKLjfXtP5eetq/giFy5RTYxCmwQmaIq
W1HyPOjn66lrzWZ54jSyxAeUvKS5ZHNkAX8cg/owtGuaCPAhF/+ZB5fFsa+6FJPJ
OL9Lu8Npe2Y4g7gpxZ7Wgu+2sAZ1TSJ6vpvnXCqui4BwGXKzeM7xjhh7wOIjiTnF
5XqriTQofX+1J6r1AIwBtmtI0T8Gh5dr4mV2C0LtwYeDMYRmrVgQ3okm1D9Rmlys
nxoYQ4qsG5peVTJ7x8aQavP6AltP4UUEqCXNyHeMJwTkKoCE+Weu+aUSs4ur+DYD
x3y59Sx8Ig8VlCcbt0IK+VUY0rqptUdZzBVyVlKRT1dz9f5yMXvbcQSB7OTRAjRA
TrTVzyc6/UIH//IUHo8GeKFqYiiGX88XJxQTHVC/1Z73YZh2LSmYKc5TtxKtr9Tm
j/KIIdfYtaLqNjaI/l1EdhTjnU8c0RW4P0mtQjrMRpZa+8R5HCpnmjK4gbqO+aVe
MeTMLZcPGCc0yEcOKMWeh/JMDQ5qQmkyVfCNVI/11mhLNbdEYgtzx9T6GyusA7Ng
FaAUSBDa4t6w7YPi4XFvxmaK6Ivi/NGJp08uZFC2Krdm3+5HQ83voV5OIOH0p9i5
mNIg+fNYPh5vONF2lupJJkaqwjBhHFiKFzLNFbm9ADMYbnAQK1+s9SGXUgQaOqnE
IPaKE2xVgFijEF3BWiEeS1L/U8a7lMN/NeZfnUopBc2jQflMbEcaAlVbMhBYgGKa
vmGfW9X8nOEbz+fiHZwcty9bPvE9By7wTTD1wb710b8PE2uwPz20hkPCPBdPQRXm
HdYTz94etmxMxv9LLddy4qb8voN1SCiA/yyWCNfkvy4ELNJaA8svVbCMh9gOuzuF
w/ytXwOvgMrHE1Na0U7nC0/XGbTz8arN7Y0qbgvE7ZU3QJ5sFqz5WDnvs9Chm+RA
ody3s8ae+9Q2fSrQg6sTdEVv/LLV/0ITTJeTQIFsJAcGQEFxRPvqhpi+POtFWBj8
psqsT6VuY3ATKhh38cBG38toQN5eivLBkVdDjFIbNMD+v9hHbOoFtFxoE7cIztwL
8F84gC+6W5UIutDqDUoZ7Ns9Q/Pi8fBsGl8sb/iwS6glgmHDSEQrMTRZv/2IcrVc
9BR0TPQ/WoaB3S9zkusWHFk1rNSxE2L4boaYczCzHb8CmpyhGbzdFSCP1SU0P4Fe
e7HIGXsj7F7/hGLIs/8db5pAKF8arkcWuJ0NGI1qk5nnGfX/XxuOm5JUh2woX9/u
B9PmVOYIuy1TdAGGwo0eiCjaRxfT6vnL/4KKTejMLIjngab5Hmf+tJD3cLGlPltO
wjiiCVzuCTor4sTrSvItLS5Z2QZngDIZuE+DLXvlPI4K8SmA6Wy+sLa195t1GSMb
aRbO6r1tvtVaW7nZB90TOUgoi3ilJr7Yy+Zsk0/3rLchLm46l2usOhRmfLQjClqL
UL+jM5HnTt1K649vgMaHAkUu8Uhk6E6uqLUxadCM246QbYPD+GXkB46DVvT5oUgN
qhMBDmxJ2OQEYxFytdUJ8qoXP3qMAY2LKRqgc5dziGyOFTFZNFBZFo6B8rKW7Y9S
HrYlknL5RFpUp3VFx/IBXLDDbLo+2Zru5tzA11/abJXIsxCSst2qEbMYae+ArSHu
kkeo6FNV7cCiP9WZNPZ2W7IMtMquNHwMk+nolmpjuJaJRyWKNxP20LOBVyQSJMzk
W82y56p9nTiKyZq2oZ/mUNuGsDxGd7rC3iaqu9ClktSTZMRwxL/8pg+hzJJ+1bw3
6XPrmCXxJOxf6Ig8OmeJRIKuaC3+EEjYiZMqwKgv0nnmH6iqKnt0Fh4YsZFzFiRk
FCtapFCvz9TF2pZqQZmhK6SvOfStH++6EBtjmuU8rDJoWOfIovt5Mzu5haXSfXuW
4pHCwcnYzPEx293FGNqkMeWVCb3JAZhAcujVa/KwCMcvyrH3yypa/zB9MEeCrRH0
Cr5ybbzshSnJd45kAcX6WTKHNKKK05fAJp7E/7CrTIgbRlkTTL7y50fmxIZmqBAo
KRnZZ+mH3DB+BOW6uICN04qZk+ruJ1X/xY7bk4WhydRiS6MvCuyzJwBqlPa2zEIn
zBKMW2TK8mQbIBE82of0w1LHopsMhxWgIJMVepNSFFnHY0fxbpvN0e29rFWuj+82
VBQo+VkRzcbek4sicGbL40Y7fFUhUr6AQmu1SH5Mv7IPbjA+MBBce/P9LCiI4ZYi
mwWVoF175o3B29Ibv31qS8aauLnc5Kdu1cBEcUBc/nvbnjOKZoNgiFQbYjUtLcrB
tDW8A+bqGnLtdknMUfkt0yuDfAz5aZ+vnnxNRU+eDwsH9GypCNRt2yFMOTNiLOUl
8ipn08uX+zYCSQTuVGiT78+4Oh7bPf2E4bN2jDsTb1g9+lLDwbwgTPH2IoW++AJY
XFzwjH4/lSdveduZFRx7TS4t352zBi0LSj+H92x+70XGBthsaVLWnPf7+vGLTKrE
5PxLS9oRFH1vPlve4cFYqYaop5qJOTvOpG1DY86c7Qx6bA1jxEJ85nFF2yNyebdU
9YJ81VYD/Now2ECZv5sj/mAyyyIahewCxWNK54pfYUYeU/s0Ov7vf0KPCqQkOG1s
YAijQJHbAoRrrs9n/5+jkyCjQZ46hvxuXw2gOWIN/gNRW7z7ZqY0lR6rX0si7gX+
Uu/D+4TNwbqb0TjFpuE6zpxMxl321CB39o7Ibe1y0zP/rf5XZmPt79Gqh62Vxok1
WI3Uz6tNELQqQB4tCFG65vCpwrwTtf9UpYlDuMeT99hbIE8EDueuK/o4hmX+fIJy
znakZS+l4PFbeWxQSB/m39W6XI+/U3L7rK/Q8KeegA7IFmkwhMb8gHeJClPc7UQ1
FIQBtwMpsF4xshCxj1a7k0YK3aUWCHy1BRcILFdOxbFkLQBuXKbbT5iCCGE1R9ek
wwcsw9sGv+oZ5/mYHkZ0JrWa58bnhuWc4zqnknXWU+Qlk7bocMaK/x55RVueTAuT
Stm5zLTujI+2RC52KFehaa5/wGxNCJuZWlO6r7u/Mod0i12F7fYUsR3VO1roR8tD
b+W0yJZjhhvPPG79r75mJ69JsXLhM6fRHj4XoKWiwbPt5/XKhYehL/ySO2Ie/hto
U5KpT5Lcc8kpfFNbuZ1YAQ6aOaGXEFZ5r2lnQhwQzhE1HOndl8CVVnWUwY56OQUg
Rpa0KPyuYJuImVnVaPq6oWPJx5Y1djlr3PqdQCftSb/xXsDwM+VMK26IBxbfJVvs
00+n8H6wan3M7mTjpaEcu3ch0dt618jK133pD1noOe957C3BytsKb0BtsSwzMgsZ
RFurOMd4Xs4X1e1VYA8va3JaDkJwMsPWeN14vvPsU6nS6S1kJ2QbvNcDGvPyGoes
w8vP/O50viMVa0+iZ7NSNhdeZ/mKnh2TMchAbH47LYCa4rO3v3QVgiNm5yWexU4g
GAkLLoK1ZMAD7z1RCDKCq5dhTyI+bbqPN81wX8QUzClmszLZzVHC2S4DYyz73778
akbyK3qjBOtFZ/la9opOWXi6/6ahD5gR7bCU/KhGEm3YeSMk03fL79DbY316yH7C
AdtOL43VwXKN1chpq1davFlsFqolNNGxvtB3HF1qSe9+CsucuZm51GqlQaIk2KEq
Z5dkOcHspPNFy2xHBxnspeXMLhcT9IkbY219hrNRq1nUF2o5TzBC+n9F3iFVv5yG
1ySzsaq+BBmuyJLr4mjDAuTRDTnS+IF6XD+fhT/P5apIZ8QwkIF5s09rDWwXz7dq
SUwJf4rE+fuVdHgwj6Meo7kTgLP7Kp8TNY/YWxsX/iAtj2YdL0UZ87frFNNQ7p1I
QQgfVgFz3Qbn0yzVzyjrrCToYGE9HKuiIvPo0OsC1K/NbmB/r7EYXmUilEFq7/4G
SySA470ordoadltybHjpKsIOXyWnj5iYLGI0FjKGtAeqHsff3fjZVwsGL2Ig6NSO
UDZsxImG6SVkvAcA776LFBtyXcykt5wR/QJ7+BMuD2nPMcf9X68/Ln54SnbWaK29
wyANPUKqIRC8YEce9Q6VAcQVVdTBbk0UZ9aW0PSTRnp90I9HlKVqd8LBHdMMGUxt
kjTpwk1X0625ol8m1FNdCSWp4aRCbraS5xPnSFlxYyB2MSLozyM9dKiEGFddTjVb
mZhO4+AsChn1WfMZ61N1u3D51FIH3SskI4THDYwMLdy9NjA+CymPs1ylcgVErnjE
mbVb/6Ornd+wHl8g688UQjGM2TKX9N+pTPm7IvlTdatH9d98lIBq9A14cah9UD0s
ZmGk7I1WJeNBJ5bRR/986FNcoRSQE/JMSJStagT8j9tVSHmkAB43LMinqAuva5bX
sOlF/xA7og2nFIN7MKQsILP9mkY86yEyNObh5yQqzAinOzfD0j4uc2Ecozqt1vae
24RtaAjtVkXbLTGC+hWdhTru5BZvz3A+3pgawbuCcXr85K1nMWZhGDoZlSNeD7XR
vscke6FMVxGugf+mcsJ4bPFDsPrTgvpDd4+/jVbCTwCy3tzHuUm7gdgY3qkE0+7J
lNAmBYre3gupXy8hmY1oCVWSdvLLdmP0uYt3QQmnxoN/1JuJNrxbvrrcCh5TdcOJ
1+GmvIMu74wGU+DlKzai8BwZpoaCvLXv21K/pRE0HSZSN87GJhvYfRe+L/d33fRR
Pry0iaTZeslJ7ETj2oYmWD2oBIiOYb1mnnWkbR5AUcw3IN9NVvt+WZWtg6Ta+dSl
c5OK+6t0qIBkv6H+HABq8NTUZh1JPSVpWT9sxS7x8tT7m7n2pliTih4SHpfkDXfa
5pqWyBZcz2SOqS3wvzP1LeaG1r6E83mWHKSJnV0z/bexWRnH+qY3NBTD7WPU+LlS
qxlzd+TF/eHrqfkNEm2VKHUjdfk715yi2GWQxYuBRBCX0Fs1p9FZ/UgGei16ixwq
2fOJ7YP8bYJwP5HWqz8FhFO9wsKM1WzIUZkagAGIcN/eZ7sBiN93roNlP9E/FM+C
wvfrQIk4JeyCMmVxRvxmmWH0izhAtQEFPPx+BNM90FWsfOmCec3GdvWavoI67GV/
61FYGzLz2LMi+VWQGSoyZ16+IxRo+3Dv+M3ag3vnjOGWffX6OZ38RUhoqO+Ts9if
WGRcf3CJNfdQCg4g3Bzywq4PnTKo1ZMb4ixjeaDzkERtBClwNOALXdXG6+xxGLMc
4bIq7YZ8PO4pknuNPtfECCzqBefpDxIP/mHByFwZd5N9bhYhT04uLWvzwhSkiZ7A
5Td6rhlLLSx4l4qKXC8GgxKauD985FSsOW3inmCV/VkhOm35YJDn7WGZE2mxN20j
gX5dx3BpcFqxvGMfLe5gkU/pWUD0qj5UaNMSpX+JQl8cXgvLHilYfB3hBIK+IrgC
oKwb1GHbBS+WdhSORFd79fYoP64sjkHaWMV3NjzKkeTo83YnzZWZ4dZbL49bjpys
I0K7DaLEDQEfhKtrtL5oGU6yh3JzFed8zkj7cNb6aMDChODJXRBz7O1C7aglgnkJ
Ih2J03jRla5+3GPtBX/tLF+ZOJIUh0uYlpdEvjk9TwsEgUg5VCTkAglX7kTk9Brr
NJgWt1TTdD904RXT+km5kMn5kPL64+yZPOzouKL/gXcxaeKD+C4jh7bz5brDkfXs
qXM+17Xhg3YZm5PB6c/CfKkfT/goze7tQ4ygLysE+gbWPMPA+ky+W15fWggKADjo
Jow+9GZ2dv0HWx5nju0yymtPdB+LBuCZAwM8PVPvENChp0134CDs5AhH32BQG1Ck
NcqSGE3iCqpGngeBloChx92SHe/GEafKfRPAHxq7RXy/NMZuNqLPUG497rNT5GoT
DcZdffLyEKyrk1FcigMZebEWyHYeYVjAxOT9XFgX3GpG1xR3aQOn0EdKP0MlOutA
NHMsX2LwG91UcESxivMscRCHLu6jK8uLXVRZUnuXrTFNxxYy4UPPE1Zsxx4XLWLz
EvhcM1tL15mG0vD/7RDn1mKjN5ytnsOs0CRwjqLO/mtjWvl/LBsvufqLmZChKY7z
ZHRgxY0zqmP0B3+yUYdyG5s0RjJZJrAO37tXhNN2RfEQGJiciZ4lw9+/SuugmyX1
2PSDVX/j7o1MOWqqjOMiRB2If9o/Aa4gjSaomnpv/vNPcKLKuQKRpVLJuzXrDA5J
B2Q6ojwyYF9YVASCU5fMGDzdkbzdZAJoMgZ+piJnX5nfyr9/e4wDCTrG5kRxU5N8
BNJspibVENyY8jTQ/TxuN4LlXkoPix/KDLm5RfZLHjch5H5BFq3r8Wf9g8uPJWIa
zacRXnLveWpfQlym+iW6xqsPkKCbJP81QE7Es/VD7KIxA/aPH0RU+TMSMhENQHPk
ZdaQnOXt5vlQfzK7irVRjX+jW9x8NaDQZsyX4p/U0Vm6D722ZtkYJNdN2UheDxrO
RHGXNHSaXQCRVIYVaG238gGzmVMCgb3wklJ415OPPkYRA+gqzN/w1CAbKOQrfvwd
CmHGY+aDmA8EzWpeiRXNm9zt5J1rSxg04xzIpmePBzZ7Wr36aWyM/6fF5qLHE9aB
KC+2tIih4lGrQTI5BdU1GifUwSdJo32g3ad3/YK54PHPi9jyMe2HdNg3oaUB98yW
pa7pUWnYgMitqF6P9OB4Gjs8gekTfMd/Q2kYeMOwjBZ/54iLQXLbT9Ty+Y23hzp7
6VXpdM3Tk9O8GCRJNmij2tEtiUSQ3le+6u6xH4y4tWf7RSNcahpLuU549ORgLmdE
ncHMntjn2PGNmrx1Wx0Ppf5VWuekvSlw0HR/MJE5taSEGfLdWAc2IvilXE7sFzD3
B2MFE49xHNbGb4sY1ZNmP4hlsW+q8TmkruuVa8sUHhi9jQAr+ZDxPHsCA6U1twJc
oMXCTMA3xBs2HjzAr0JJQeb52SRaE6OpqyozQVJIpZDNQwSYf/4Ph+B4lpb2S5XT
HyUBP5RtpCH5yK2pIdEbz7/j3kuk68bX3sVQeQi7E0/mchr2iPyelFAuTJltTpar
VX7NX8d8D4HD9mWs26Vt7tG010NwJ0McOMrDYDVeQDOi8xkpFE/TsNj63uGu6I2d
+Qgv8fhLn6DIXEhJ8DPWYz9Pmw+3m7oc3GjKmjfJ/xPfBB/+hYAxIUtpzokn0NRc
7KG4Wz3eW3wBXFJyvJ7E/bH3+YZuvsZdVIizDX3/WCfxN6SeIOdEbr+wgqWRwta5
14CVEQ5zVh2wcOIW9L3zTbUkgh8Hp0ZHw8kYQplkaXSr6gRtsfytrSctvnyCFCmC
VfPrSQiTpqyfaIYvhPWhn2mLFV9xeQmQTk9wNo/vQjiyB+SzaSmFoOhpWzhcy6Ul
ZD2CJxrz4KtnnTcZ2NAyS9eMTV+cwqs3umBu+RyD07WrEOV4u9hdIU2839nesfMZ
rLgXIhFtAfCuO/H2RKlhsyFmJNiOm7Yt/hQD/XFNEC4Ov9HrQ28kQIT8peA17Wyz
gjqWBPotin/5FUFptzfaUKgKyu1qIKa0Uga0TZi0SPz1jN/lDGiOPW4otmaj8H9S
WupFJndUFPhtmLgSKY+nAUDNCjfig8voSSmFBoj0JaMjW1P8KVXEIojVz68Z8Bes
NEzl/j77iPEYMkSnm9tDV1NMKQKicRnhYKFgSbmUdKL1QQpWkxqEzYyED9Nj8qcS
3svFwJFyo9WuymH4o2in4MGJru85trq72VxNAo+czMsMdD9Qghl/mf/jMjw124Ig
ns9EICPp+vL1gNEXZEJ1KQhAyYxYoTdZgIxVMh6wBagB9c4cOCacy9nX6q0jqa1f
4OTCt6LfTbx2ALFFxpJFNwMHpOjE1zrRku9PPKftY1MBlVLQFl5kS+BYJCGDkvnQ
aRsZSeLLMmj3qEYLoaR7+cOfLgcRGw13a7RIVu9rpOY6sPMkiqi040AJphzBjBmz
kAXiHOTkr564LsDU9vW6hUxA9Y/PeLgyEKNlxjznQwuSJ3DGDDo+N4wt44JSB2C7
F+AVLijoSANCZTkcD1MB416WWx4o0EHnOoxbTKRn5t1qYW27GKHHbbYmbuSeJKoW
3Wfc/cbxFZ0DpjpQj3kQCXNAmsUOsE0jjN14RPQorf7OayfK3QlwDPtfRPtiiRq/
TuF0InK1t2Ewfd3IFAk8ql5V9w1J8qDzfUYaRiH0sEvf/Lyv/bzKdrXCjqk5Yunr
WSg6jo5WkaUjZlPhzl/kKVXCYEHUIhuQZMISRM7vi7vPHFOmwndr8mOd1sjwOuZf
lifEje6k4t4uWF74afyHLgwQSivA4vDz8JgeL52zW6T26MmUzb1NSZjw+irpk2GW
Z3Q0fBmirRjnLn+VMJ2uz3Qn8e1puc8L2s+k0HjwCNzVYaBATfHE7qZcJ5WH8m8/
qq7TWyYF+j9omIDwHERNoEq0mMjKo5EO9os/xV3IMsPYwFi4HztMxzLIwB+ZhDhj
nhB73QHV9jRo2eVhmeRIdfXLXxSzqO3bcqaPrDgYD6a79DKvINuTF0uoEdRVf22q
anKNxg2Vz5lhm6TSn7Ae30JNvZF7VcuGT4cAxubYhlyakaXccu6oUH4Y8bAKss55
ZKYs111UGsXlueTvR+miZSG0HAngx/EYi8g7b7u4UJExsF+C0/zx1jgsbqSPclA8
ah3maiBR4mM5aDzjAemgyuyyTJGjWyq1SSVSg/WqM+akG1KRNB66DnANCvXVNeh8
gafLJIanG2Nh+5VpE/LUMGwl0IPNLDBHFuKx+1sirDykR1A2MpS2KAT0Nx4hBFCb
dCvU6cqM9CbBWzfBh+whBA+G3gPbl9r+kUjcwnYHiZfwL95e4yPf0TIdM+58Lypn
YhF8a7KsuNiJDeVbn24XppphL09EmNIQMtG+ZWtFWvWDDDP21mjMRiLz6p9YrzeL
IdPQtWGmKyAzNZetT68C5PIZh2zq5JINiU6OOdM6+QfjqdVs8Q0I/LjEDn+xw6gO
YoZ70XINVrhhz1Z5qr0ZxfVm65tevU66xxaR8ZQnvj6ZQBMu238ntG1t43s36ygj
00CH8v+/GN3QhXGZJ9B5XaA6vWBkJDhB+CIKZfxpzv5/a4EnQ852x0rrCkpHYBoM
0p1HyZxpFJ+gSb/DJrFlxZqL+oVSw/YhtN6YSMk7Kop8jUohvPSz/crNlGD5+hWh
hOpyprN4F2hXcbp1h+u8/swqYPEEuY4MCWPHGV0SqIAdPNT+4H3qXAaPvKC/pZDs
s8j4uNDMweoH3D3FspQU8tOFyhz4vuploxPG3cwA2q2u3x3KRF3ijiIeyWgJLmdn
jBYh4S48caaOANAWEHg9TmvsHxGvBJZNSWtZrK3oM3SalqMMfXRBGX2KRV48p7Gl
fwG158I1RW637uIB9a6VyBETYjgnMQTUSxIg9sxALpceQRkcRa5zmsEvfkHlhWRS
MveLHxXVBbiRcvm7/ffCnCjohE2e0TTGKycR0KJaOADqcmQEnt158sWyB38CalHB
jCYptS1pUHXzZAJhjDJKoQbai1qXj4gr1eZmbE3MnLHEEMYPdnB5WHuAZxo8QIfO
YhQxjwzqULN8AbcR5tJ+CATiyuzUvf8BLLKN3qwPOTyeaIKlsENk0+I/UrJolCC/
J9HiSBX1aDMGKo42/6Gf77g00CSSD3b+2YZGyOwE+xUhz547yviE0jk4lvAF60Ia
Ffa8CFoEFBe+0L8xCCtpnFaDPNwU96KbPvT0TzJhifRaXThlP3Ho9LuHduv/nLGa
iCTuzRBMRE9PmbmK7g7FE+3IpwIfAvfyDRpTmDQ4KT5ZL/WTdlJ164DDWBWKySTW
9q76Dy0A1xoPCULz3Ch5yAToEevgyh7RLUhtvTkHT0fa98a3gyJ/3Mn04Am8MFAR
kUYXcL+5Klr5Kr0AFMPvQj5vt8oqnzz0nOOSYvrQlZhkoaYR8G2PzFY3T8saneKA
a+yH5wfjY8hFtgHlpspmfoe5C99pBsyrKn+8FLc5JLh8gFzgv2ihGR91Hf0/m/bM
njCFu2wXnGXMPpoxRK0ELB6dcodXbIQQjSJPLHBaWxHVwfZCRvuF8az+BYmZ0u1Z
IkiYOEN+2Qe/tktHFG2qSDqBiF6hPTLfON9l23lOCOvAt3BtMYpwodQD6eDEskC/
HLQm2K1auRGlfb9bcPjWP0r797GWL0doOhTdFWRgcDcSoqC0gRzbXcIy026lmXSU
Ewjc4XPHcUz6RE8yRCN0tbrk/pEXloH8DZynhypmUD5NOKqOexY5GrKdz+WwXcfV
DhEivlGQR2KiNbeIJtf8PVGuLo1mVELKpjA1EHgb0c2l7Rx7+q0g3/S4VDlMdFUC
CmnmqYPwY4pVVUqY85IvmXaOCSFPPhhT8n3mbqwCtv3cwIrSeP68M2Kr3QXaqzca
OMdNt9sU4NrPP3yWpF4AGWtNE1MiWE0LvnY5svgC1oTWjkWkYfUKC/jO68Thx0+/
CXFv72ub4E088HqT2FfWp7lWD9J9T47VEf1TMOjYQFMBRuYyqjE8yoZVGeoe/zk/
+2MJl5bxTSsOO7S409IOBhBhdOOyaFXCz2wL3Qd6r7szRCar6S+leVfc34epncuZ
JtqfIQ06E4BWcnDoBAhkWIgpBXNn+59vvCJG0U8h2wwJjYYRqPPXkzMY/adG3bnB
yieJjIkNwZdsNjFHNfFJY7+UPmdosnTMEOEeRzSkhSMAKnSV0/klSL5IQniASFuO
vFgPZxEqNJPUtwH8qvO4iYSEtJdLPvCJ+GiuW9HtEcLWsbckOzCnO/BJcgu1FvkK
Ag3vsLXWjpHdn3aWDR6TfxHCGb2HKhUCCYuzY6aEoNGHAAvGMOYCaDJdK6JgcJpW
ORZmK87Sf4FmaSaAGoDe5SqTpTg69S74vYwMYaHnhVf6IUK7reUZ0Az5XLsBSJVl
PgMEzveiDmeUgtVgZpZv66dd9Pi2D2YLU+qfiWMqUh65nvNkrGTdUUvGt8UQtJZ7
JWms+dGphPw9KuYg4Pp2lYkIlJydd+gKO7QF5DUN4430/GFmuzuP3gkcxquTTMKm
cV8Ree1Cx7Jn8x98NTSrDvXcttwbnT8crt0k9RHqHG4ZBzckPH5r83mpoTypPMYt
v2BaopIQloFf9Fow08hq795209IOpHWFqsgeVkzLyx8pUTYAu0nALNb5uJMfP2wP
C4ka9CWrag84EQxRdUEAp/1O/SYzyZ3Zj4yEZvdhb7GjuZeDGDXPz7oNZaDbaDPd
5Hgt6UOnRABigciIZXo3hZMZTeR5u4XNQiDJ0Q0n50moSmbpy6vbgDb6I8IuEXx5
I8qLLg0y5rmTAe2T4LVMzDLi0w/9BZ781td90rOgIeOHDLNHxfqdQeScSXboqP9h
unKWCi8itQIfZaajOdEyUcF3KP3NyUBin09e7dtCx2yom6qmEpbx8SkBIyQjdCK2
SLRmhe9M2UJRt+pwYvD+ReQzTutJVz9EPSqIrO0rxGh9jG/0d/cjaoIFgtubGzNt
odQixn+xs0qnBVL0MOXCx8aJXLHYv4TuPSkfdzIKV2YH870F7INVFTAJ5WZA81+F
y1k7yaS8NjAIsPFkMMUBJPAXyt2BIHogV00+2p+x8snidhuDdzFXoXN3BPS3UyM3
PrylgpoeKrSh5vJv5YqCeQC4U2digd6zyAxxWZ4TabajLh6cqqpF7nkNEwM9svVx
77MhllWsX5lP2EHqm9JHIWypmmBsA8ci6AffqioNlme4Ndgmg/CXNXlMhh9Nds2N
/sUPN4pXw5R93e3VdoKEgbTxHrYkMJDFsE29dx5/sxN+OJee0sDGQVDat5+4sN5H
udYZdai5J3xgV90k9e0OgD9OFOiQoYUR9Y91iQ978pRHva84NyLW4ZgzowoMIDBM
eqhY4fcbYSnf8oEFRpZnjLfKvcD3iEZseaU604A00Nklrr1vsAt9gVkNxt6PgENi
mZfrylJBHfldHjCZJzEQ4gRYW3OG45h6QcdUvnfE4BQEDpZ22CBU/4H/hnpT2InJ
AcvcD28XT/OmTmNh6EGXb/Qgaf/3uJSG5U2ABcNkRAEtsFhmVdTrcxSFNFZbJiuh
Dso1iS5OQRg4rTny0jnSZFFARezTADwl8S7A4Q6auTFC/EZ0Dz5PVigoZBIS3ZNS
znOk3Jr/j73wCvPPXefPn0vial/WzEfwQ8AvclXC2xbKB2Jty7yLwL1989roZwnm
ULApP6uacy/knVJvHKkpLOZB6viGPOthmIb4cAQk+BEO6tmn/QqwsFOUJvYN/jDG
Q5e3L+f6o4YNUbERaNNHIwwi4Z1Ww5FCZPIBsKVwVCo1bEENqZE4LAsufYQpP2vx
DjP8yJBFRSaFm8z2KKxwEKDcnCIUnyj7JaKOXopQDgLwczAKszVN37NNcHFZ+5zd
Jec6ZAInNMIaLPywLwcNM8zNx6tsrAE0WsuqQTYRHiNPvGunjm16bgWivLUTdXGC
3lR/iZ40a/Ub4zGHqxwLPQ2fOw2WTp3n8MxohGiYEGRLTeeXaHeD07fNXvVTxOE2
RnGKXASbTkGYSQto9BdHB+9mJAwsPBLgkTwCVABBDmlT6RWkmj+nTjCbtIelnQ4t
IaUjdDUsQs26Tz3lx44a/NIMJMpINBdK32W4mdYDonjjejJeqBV08MYaEuaT5a02
Qfy+8czntz7Tfwwj+QDAx3q4//Szui2NdPcDTEXs1D4byLyaYbE3S56EVLbrQGTf
ohaSSkDVtP+nnUX0aM83utocUM+QGJiPunjDIe8HF0wSObOYYii9UGZtarvvqXqF
/kiH8haUT5q3TvNx8Diskor8Q4+sMBHkkv7w04J1AsA6wJoglnAbioghL5fzXK/u
P7gZPk7JBefB0WbT6LL5KvtwCCyOMwFFpAnACZLtycFdrC2po8Osj4kz+G2cddrz
yMTNBs74z5Azfyw0a3MuQ0j5Qq8fHT4+r5a9o8XDidrS+1HySZt6grjqpI+HhuhX
Wfu3eTPBgyYqACWsW3cWwqRF6lAp/izSiW8gSRuvvy6e2sIwEZ+BrsBF6W4W867R
FxJy327WZe2gpmaq6yHnvP9g1vkyXTFZY2OvM7WJhnTIK8zK0Yjr6EczWFewDkE+
8sTkIIWI4J6i1m7Bpi73kWsX2kpz/WD/HJSNHiFMU9Rg1OyQwWRl1lvR4B1r9coS
E7hZXGfwyA44e7UOYbvMnmVzBosx8oxK69t4XlxQBi/X9CKiG2Tn6h5vq8rZzy7K
ysdZ+oTx1M6VoDKFRhfdv1X93Dt9CkZOW8VPqkuLlR/YjRSsbGJjEtLhC/O+WV7T
s2GUl27yi9ymOx4m6DNdOU7y2HknJ0/4SrF6Nw213knyHZ34hyJ1oY+cXWsoiWkn
JWlvY4gYJuPHAr6sKd+ex6PkWVA+rPloSk3N2LYniBLLU5LnSyVQzbuLCuGr8Hrk
dE3D4QRA2cfOlsB4VjjTjRbdsnDeQPjfq5nbXOEvatsgIiHorapMHxNsC4zuCQ6i
fhJDTLQFA64SpSTPwyaHPrN7mQZ7gC4IjyhBlUBytLql6lht8h3xABff5imlmYvy
Zz/25syd4QBKiAhSllGYsZJx1P94e8pfbjyvV/blV7YhTf5w7yVODHPttRWyxOVS
WX54e/LSReDKSZb12VbX7YJMWt4/wM3gU+DLAG20dOTZXaAQKvgj2nAuWpkBhrel
0VxezAhXgM/u9t2aJ+Lvaabjjk6Jy6whAKBa22wQyVPmn0a0f6QDstOHZ45s8YKq
zMET0WnoUE1Ceq1lMoyTsdW1ZbCmru86aBNotVwrkJ9kvFaZYh/p8OL+ka1RK9q1
a2+12QHLb8LPVI0pFBMafAkutrxlK+s66MvNgdA57RqY7Ur+2rr3f9PipyVmZCL8
/zj4UmNSwZQTnj1Hu9xSDAbWEc2/tMT0xnHt6j2KBBuBNbj5HWYyYOfKia6U4fGW
3FcDmjSHcz4bZB7mz09i11uWAFisCs2yIM0jsq7/esQ0FqI3AEBZnezemnbA37Af
t+qPTHIcy/SCRBx1Q/dKwBLJVzfl9jGLnCym7K22DVCA46ApGGEvoMD1yt1p0U0k
6duvkqH6LqqFJidrqcwXHQD6741TNEsDIvG/Mcb48E6O9Efte2F/y1zpH/krBIMs
jfndKobh1WdHXZE4EB3QKZ3DtRPcID7wCDQZmdftIJozjP7BrH57s0H+GM2xhZSr
tFk6O4R7gaQaa8FxGUIT9Wkow8iLIrB1Hy2naQhWo0tsySoNexsl+9edjCnPkPjT
SyC3R8rG02hKkWEUTCDDMRLt7zhpETX5Ti15q+9lLeq/UoFGOpOjQR2POG67WfDd
EZWg9MLxs2WvyFBwwRkc22pq8Vl89l2BzpbQuDEXKz50hV9S+NzAc6Y4l4opFt1Z
HtvAYTAuvVnlw/sTOWiTXIdNsquTz7CECHKMDsh2nJqiFqtH1gjJI9H0vvINuC9i
ikv+eK+UeJJQ+UCdQXWglVJTt+2fKqwXJ5P96CfTaXlsFgyRjHHX1qEZAVpmh19y
RLLBQZhEm4/IGu/BoNtrYvBgmiboVeLfYCUL7AVI5j7PpwiXciM/MNB7zjLedmyL
1CmMTJV6MEpnpnTrE/0gMZjuCwloffSjpm8sEzcgkDj6ZNE5pcaOk5Z0i2Q/EnHx
TSXcsv3RBxt19MvrW3if2dgRi76T0wdl94XizYoFt+bF7QxG4QqPX0KFFVDxEZB2
luDAiCU/e2+psFEVqsGdKFuAi5HkfmIxn+wqseREysHXbf3OVvT2ynW+Kjzc6H2m
SNFNSjU4OwXvhUnwXffdl/WgwnYcSDY1ElCdvNlSGH3BoFtqsbm24aBhwQjYF+Ip
G886U/+kDi9SwgUSqxGe6OtP64bC3HHCmsKl4zj9Ma3hVH9SyT5xlFMh45NYZL5D
7buwQW7wuO2bQuy146fFlqreEIhBrSCF0KKAFdV5M/INUzWtf/3gbR7BqXW2zbln
fRWqyA5aYJywZwgZr5AaUO3UahJeXJ8QXSm8xLi5v9+f+P/AYMehmiK2YOppsmTR
GZgQgjtJZSBc2z7aH9fiFPoosbkxFW8tKenhHzVzNnZlQuwdtJIoLGpsTEQfj0Ly
DJnmrKjBcoJ0QjwaaNakEfA2Me4vQWqW/clvmRL9SUwPeTg7QjcdqP59iSRqdXl6
q07QFCiHJZ/k5pHWvB99h0u/b8zsbz06QUOOYXcAUZbAEMRPuYTWURiVfqRVrPbC
lGtbjeCOkReCGc4Izn0gYMXPEIEwIAYjx+c2CGdEwtDotDmNR27LKjF4m5Em1YrS
b7xISk6iDlqC4jvNW2LwrDFdQIl0GU0mTzI8oCUaSqJWNa1XJ2a1K+6YTHf5F2L6
QACc2jO0KhRrNwxRh7dXOBOh1bvXu5f5/ctQc+PEKpRrwcFbJMyS3m56CRdx41yr
Qg40yhDgQYRPR4iaImbGIPRSz5G6NJPTYxvowmd16lxAWN8LLPPOG0iMqMKIeJye
4/ygpjzG2pjFvmVYuTI5CMExpM+uuo2z1h7pqL1BggY3xH88jVAUPbXHFf1WntAR
aNc8f0HsMx3cIO5htXCR+Zd2PayQ/ig5JyLpcUWVgCnZ9WFx7X6PGAMyKWduYv8X
F8U00VhRISis75Qv1nbFbmYYYpiAolU9y0mgZ4obHYS1OUQgi/wI+1HMnviY2J30
Ta9EvUb973zVbHuMbMlHR4C/XvGcbYPBX73zwVZ6rzdqOhFTEkHxMQFjoPnlcoJK
RRU0eyhDeNRxIH/ihNnih/moYThKvKu/Ikpnyt+7K3qm8b0wtSHhjyquQJdtQjKr
oBGXMFSPBxzYsv6XKED0vnWXqBA4QKqxXgW0z26VyoCtCwj6NI94sUlAhXXuqE4x
l+s8YRDbYFSUA0Kagq2saVVR50ThmaiP3YwKy5LdS3Mzoyjym09td60YcaOkPTNY
5aYpKtaa2lrdJIfMzUbHWdx80x84OQUiIromL2lWdrweRSc2g3g0SUtjkBAi4iX9
7fbydtU/dKrE4GyK7FESnmOQ/JXcy2mfcvRaciea2NptySwrvW/S7qioWd70D9Tu
nkMNMERU6s42vvYdOZGpASDyDRQDbRkNBWa3pLj2DGBESxX+jfEsGll9td4mQWHM
YzFkUe7WQ672BPjEgJD6K0dO774SF/0wHGiaOCLqKByrhIL6ljDI1ljBOxWDDT9s
WrLHHEBgxwIB7819qT5qEFh8ojsk0yQIlPhFa9m6pnEAd5krBiWiWDSNGYQwg6jU
1eiDp52UUuc138q4nnhCKHHvSfPz7NH4UWyTLO5dmmu4QM1v8eAwcK1bxjcOwWdT
vZJ0cWOkpnCSRyVbXbFR5enEu9eGX56ZqIWiLaKs/URvChAcn5x/Iy3RThFuz6Al
LR9dpe0EKoKdZamfRFiFLXspZ95Tj9GuhzgI6oHFOPbCXQr2op/iV5mgcpmaHbSr
XzgwBWWU71RGxoxrRXJylmjrx54ehTzxFhdynbTlZJH8FeF1GC8lUgiY2WnpCKMB
Rqc+jlqXkGlXynOtqvb/coxdTy/R2aZ/bWAgJ1srqQuXQmZIaXWhzLkj97tzPHeN
N4uqX0yen5iAD5FyWmSmDoG8i7fguVa7T8J7006UECcThv0sRssFgZQfCB+OPm1I
OJ7LXA/nWMYPT7Cr5twxXbioCrHbKfu++miuoi1PVSBch3PCpQG9WlcAxkLJFWGf
7WXnRwKME6VOTc+QwKc54hTEjbWM2R+M20Q0oGtI53CH5fLdI5Y9JrXlsPf1OAwv
PSr58zd6o8Ix7TPJdLFnt0QpEaAHHcM8+FncANRZoSkEOsFnxRWki2CldqrrG7S5
dutbQdLFFIquNuwXHhXlV3mbfL9LAWsnCiDN95MxbQ9UeXEw/5jIbLK21q1AS8u/
qRs9il8K8Q5lgxME0g3FIdxusqiUJHrO+V3en2nSwwvL+rQvmir7dqOp+bkf7qY5
Aso0gWikqBH0pFU9GzIQ1nYVlzEhMn8AjXAJK5OWR62KZ3pdESoO9Lh0rBw6i3i+
sIc/lXunou4nUrs26PR+wm3EcsWhXvHJUyM3i/B8a9b6vb237dnJ7nPAraBeBRMW
G6932v2YQ/Jrb7dPOTn9aO+fbEsd/U/MWGn+07w9aFMG39Wqx1RZelO/i2y2c6/O
GeeEuNdPHd/21sDS2h3uQidn4RAKmrDMQw5OQKOIr9XG2bY2Nc5xVtVNHOwXdwuJ
II849D/icrYnHTCPBZWpjAADUQDsJ2V6fCSST4bvSbJEeb6FZ5DNZ6sM0bEKvKc8
VBWmV0igYLZbA1DtLM4UbmI4obQMGsyrRClfEaKQnuPDrLxWTnWI3DDUhq/Iw3Vl
KdjEOdo9kJ6V7JkhWiGS6YSR1H/8xrFNy17fPTNbV+I0FsJADbhZbLRAk8kuoCsq
gzX7I3wM3f9OY/odvWEVEwnamoMdOUz5V5yD3FhUMzFmADuKibA21Dg4bOrCMVl6
wfEACkdJgoAtn1kio7Cpn0LN1kbfyEkxDvgcALpQScDkhP20Eptls3Rl7dZ8YJcn
vzH9wN6FIzDU1Y3/uaZneAx3FD8x2ns/Ttf3/IQS8oP+yFkLKW8qeC4QglVNufJp
KyNKXOYRJz+U3J3raX//Q2KoJz9vGe4dCvYML7ntBGPM7R1YMXtj50IbtDW1/iEZ
cLQIiJKsEGvoDRH4YYDuDT5I0kGPg3QuFLVDXollyQTtqaXGBHngUy+RuwYfEcMX
MzJpb5NmqAeDnbycxxJO6/mtJ0AfbbuWmwVLGpwMUQkpr7XP3/1EIAxTPLbuK43f
uY1GQ98BvgeCQbTbmN2OmGbqz42R3zEFF8j/oai0gnY1ZghAji/ld0WeLQI/1Qpp
cfKsLFkiMrVXqw4VWzSLmqvYQ2Kmpjzd73WVBlyR7UcQsO+G26zeHhyaJJdk2gi+
uj1LN8bMCXpQWuo5Ksgnc9A3wizDqu75gEZNwsyBXLOkjC5d69TZIJm3veTN6QpP
QfHRsN8ZagoHMvnbKfB06I3aTw7vf40xbnUp9wfP5wQhxwC75HmeQirZbFMjwRVh
Y3meRU9OjC1ToG/QZNJkyiTZSdNVwmxLFQFO0oo0Ljz9EAEOjXdYJSTS/Z+KF77F
JIuttrY2lnCKNOcmAh31t5J1uWTATZh5D3alNiAeoGx808BSQOeo0iM3Uv9rXd/i
0cgRvb6/Q+qJxp/BmmW7B3JIn7BO7QLyw92o9mNxoFiwA3RUrwYDsBrz8lQsT/xL
s0/eC3xuLb6SG46BsfB3t3lTOruqMPLAHXxEzmv/f0/5N00ynS3/JLutW0cn1Ea2
okoDKcBCvKr9y4AFpz/bywaEQfUcMJPVW5Gb07SA4RXgUiIWngj2KYEwg93YePv0
4uYsXxG0A8EIfxt8Tl9lQovDL+LI/RH55cnsiq7F4e5mJHTXTIs6y2vWoYWfBLUD
8tF+P6CRT8E2/zjAxdpiONaVG1fl9oSq/06WYV+PfESfchqxKGJkKzoOQl0zEZIi
WYg4abhojs9yvs0gY+ZBWxCwE4dvxH8+ZPTv6GXU37tW3K90xZszZosCdpfs8BeB
t7dRzXbH8D8V580fWvSbOTC9h1ErWrn1kOS6drwbszTdO3sRAjqhZ51aOd15x/xA
jhCkX1P4qwzA+FjkFdnOrhAJHe+z/Vc2K8v+kOo1FkjkR9n3qtEosbg5Um7dUupE
0egmeNFbpUpeQ6TeutVVdk9lTJ+iqVKEFh46Fn2+tMNb/zugoDq2j0D+W4jh7JzL
LUj30pEP2EO4UKeKkVcpm6gaGvmA0yeLO2OibnTYBMN2StMB95UohYmsKG44hNKS
7AQLV9uM4ZfvP9+PjeKotoIWw+xCygNhWwIUVBUnV1s0nKbJ9a0Iy6UNtn8ny2yQ
32s/ydfc5wyJDM2VYp55/HpZ9FJnQncVFBl2tVnnvqDlBVdx9qEnMUi5M1HHlET2
xP4PZ58LS49UGj9qdvyRj3fVUSjq34pXEGjA/ObFmsRl8TuusRbf31BXOaraExYJ
YzT1pPjv9q2p+rN1/P2TuXZ9nMZfG1XdYz+3aNwJwKguVg3osWcLzMpuXvdKwg1d
5B6tAvvUN40Yt25CEPIHNEgDWcax7nEfPiFJmyzMlzE0A3DvFFbZdH4USVLChd4E
LB2YX6XwxQlMsI4fEqs4eOyGz5MA2SAPgrDuuw+viULN+pIj7HSd+6+SL6L5pi+6
4g/sx2TF3omjA/+jcpCIgiDpsOHZtI1iGAvC/O5SPnZ0f06voe9nSE/jONxk/Qpb
W7sF34ouSkPCWP6sxqcMzF/PT6iLusywsWKrhweKdL67UVMHYCe3yP921HJRTBSl
/TH367MXWSMGY+GTNKs2xsQFfME/VtLH5HM3TUYXAjn8vY5Sbd5Ec8Fa05zm4ZaS
Z6ns5zW7FvL4jQXZI8DLcoBisBNWREa4qBBnLRSNTdWRtl1H+ixHTMcuhPRT41WC
qSdVyIXOkOwgpLrkXdr9Wp1Nwzfqjc7lQ/m72/9zDv12PYhqma9xKePXUkKqkUXj
nLV0MZ82DX9XkOGNd1szfsjFH62KyEqQAmSMU52YFLV68SNLN/c6hlvqQVM5v/54
NHJSHlIVcmg8Zx0BjPhxmxUZ0RrgTw/OHRCDCMqIYElMFNYSN5iL18Z228vK9qLr
OlIb44gciwH3Achm8dZl+pcEyvp5s7c1QuwUJSG1WMAcqDZWvpUD0JO/9G9XxtDC
iP6cARFpvZ3GuItLTOlv/t6KZ7d1zEkq+wFtI8wEAX/RzbarFrueMp0qqQY6pBme
ogNSEJvglSV6Swxgl1LDKWoVZBRPBFk555O0tCDMp9VKzjwGvbp9DCKRFp6+kHqf
beWUz05sAGmnrHKlheVu4SqsmiksFAxL3szgEqhTjpCks4SOL8xyvZelgGtet2H1
IfmFQ1o1y4HUv8NDaKy3kMm60kL0Z5PchusHnWFtoZZ7Rq0VRkhwh45REwGxBdQW
NiYQROnuGEJySOu05yMKQqrr7UI5WPZrmFupxyCGQqbUls5v12W64+w5v3ywLF36
xGZEk4i1BX4e9wA/DJARArYKOc4gKWfPC2nzwuHnDs3awUXZo1J4s1aHPBO8AxCb
HP/XGPX9+EXRPFyIsoSVvNm0Ry8V1PePhAWsyt3KqYZVYtWlvjWdzzkeHZUTC3vG
DpxrR9eGbYnFRdxlvOR5InYdPRjj+n0b/aDz5I68PvnO3PYbpjZQf3LpYPilzDsF
3BMvtUp/Psy4XkUO4V9CNMM8oHXoQHEvz9FmB7h0CBWbfzYB6SeNMYfBCDtrRigw
kh4iXGqxZq+VSYNLsDKrZ6gFNrm6DZo7nHjlCmn+1Q+IPT5fWezAwjXdyfVTjF9M
UyDsQbFCKXt8iJTNUANZ3oCrA+aiPkiRxlQk0FLg0cpuMVmO4CrX0649jVx0Ylca
gaP0SP8JT2CPnkKpuh1Ll5b7rF5o0+/I5ycf6NeDtzS5q0DX6RisR7AHWzIP/jE6
W0vKPQ1YfYqKpvROPN25wGKvDXL6UUWAkVGRQrqdXgiA4TSKBx2cVZuRyM+vQ8Uq
OCFbQpYEBVKzFc8Dvf6f/tkJja27uhezxRroDb+9eMRWUpamoFDeidTkFxdzmCxA
rRgjqBhpWxbZPVfFXEtHCI8rA48ac0MCaUxPJ5aJTuEKxUj3O7HLvnKaG/+xlAP6
vwHDHp3pmJYYJjx25ugysIKRTNrVp/n/nTk9903JZ5PKbDCU0FW3XHo8E1nvh05q
1sU3AwUJEAxQA0VpKg1FwvybSAt7q8RcxJa97z4L/rCB0a/Y7FSqvfEbHK2xANG2
ymt4K3hwZuZQBTJwosOjlLLE+dNqnUDnIQTwy/I6FlpwIY4Ir7zu/VphLyfsbRy4
mJDnzxiZxBSVU/JdhJeMWO9HoCF8/AyNAgTWjEnVtWIYFH4f44DNP2pIocTafe5R
4UAzS/haK/Ob9PFIrlUW4gPTYOmna1XR9KL1PQbfjBEdubZvK13/9g21Uhm7oMPC
9gkQ8eTZjgcU3ySQ0upbvcdF9XE4IsXt7IyUYlo61WSmdElsi/nrR+N37YRPzofO
liHrd8ci6lkF6ZzzIk1t4upSMY90MBFH+A+b+GGrNaWH+v91GtNrkz2yp9/RNnrl
P1TaJIMkXOKy3fFz1x90wBRqcuFbeO9Bch058FqoeVgb4bx//9+mOnwK/oEVpEZn
5BOEUX4uaLExrle2s8aKTwyVKUdr+ZUHtWCCZ5MDmRvasyINOK5FI3UATRBHl2CW
CcGN0Tl+TdpvZNzUxahjDL0XuWEzDaFZFqdx6nhQcEcUFZsm3+x6UFzZV9nvG7vH
4hKrNtmb6t6MYaFkFrtbTdThj4RR6U3CJbtj3wb9IV/6pYeLasJLXYAI1c1Fbrrq
htyhsQUHJ5+oweDxJ/zY7uW4QeT7DlMpsOYqNBXcNsMTCpU1jhuNgyHjqeMtM4ZC
aiEhwgKpRjVFWIjaPWj5S98JJ+ET7B7QRC53Ex0j7sI7595/yGXixJ2gVf+agm6l
tk+uGNODz4QTYA0DnWObfi49PoPceHF2q+ZKgqK9VGGDixS2JqLRCatJNrxnQ41H
/jESzfkJbNQKLeMjbKh+UZUl1Eitv4PGF44KWkQZysWeA8LiFDpJXE81D0gLvEFT
+C77l8Gejz1qd939BJQl/O6pANSWRJQIDt2h9OK9MGrsOSEwaE7My6NAPHFZFIn2
hImgXfLuA1g5qLmOdN9rgUXWeXA0Co5Z8NENjAXakAHNL2AiEhDLnImWv+6GGV8T
5c0VXyywDiEfLRnz/VaIEwIzgwepJDhRcyB+xyR6U/lSLMvafIjwT3bmjx/EsFUv
3SNKhPK8zMswjLwuvlo9Jfw0Hr2xu6rmLrYAPSQnK9JxsBggNtFNPgqajna2Au/Z
Lx46QVxbUpRDRGy3ICfe67snXsgdYF/Je7ZCnJn+p0hJ1poQ5YFFyht2EyTsR/kj
J/gt1AGH/3H+M3XCBkcAFFuacB7V6BhUeR3aT+TwhHcVmzInEfzTZvQV+M9yAaGx
HNpYPqseQBDFsvfhXbFNGvA7Qf4lErWOrusRfqsKjLuLSGh0PecZ90QE4pGlU1CM
s4g3lkol7plyGlofKyFjYv6ef9QCooTQP+UGeYOHYCbAthSsmUXII7LpNnaxrplU
W7IA+NJibwDtvwHfYZBRKPcCLyr03MBoJXML9A+Y4HOx7lb1s0kjDQ1hQA0lp8t1
4ji/0NaTcAuaq+zxxLd1GzCU/FjcKOpHce25aQKRdzusPgH8D5PJnR+mG6Ik4kDl
okVHSkNh1j72mjG34p+s2z5y1tKFofnKi3clzqZhudyBLJmqMqTLtnvUVFtq02Xd
ayH6R/tlgRXHVeC56DTQJUVRGjmtrxH9o5GvYVD9VHFLCkSel+7glABz5oCgvcqw
PqQk3RqSYR/G/kJVhopHKS/ReoDFdh6FkUXbBCr2WgzbWhht7lDXkIMoHdrCKH82
n1XYbtiXtfwVEZXqGraTUVClu/zJ2u8lnayYr5colmyjnTuw1wYQiDbYpGnlE6Mr
ieC6beB/ROxnO086XGGq6AP642u4auwrqcX3RoJriBIGJ/awijpD7r6loineigbG
yhxMVJ3oq2rCg6RpuT1RIBwYL1ucwd2At2myQkC3E3VrM3y7LY3q5tpWzTG/gThj
UXkb0pyydKONjOD5iepraHgaxy+49fGAy0VgkIuo2+Uuo4zsMXSsd4ByVfVcHi6J
dMSvMxJha3/SYh4MlPMMdq7CB3+/dXX7WwVN+99xNHJWRc3XC5WKf0rTwIQN1v6Y
ClB51u8Rl1pFvxpk5fAwX73XuvU4ZLVhZycO9POp0NIFD0cG4EucM8i7JvXEZCQx
atLQhHc5PnI6mxhJKwE6xkdi6VK9PgGvvpWF/QzUis8pBrdks19FUiYtn2H1NiBQ
+xBYF/1Ke2VFdzovAtToFcMhGAia4GSdPi1z1jRJBdyFJQYIi2QGHHTnl5BR5Hg/
mv6OWnCQvoN8Ww3BFsrcxQNJFTpGq9wp7idPi6kK8mI6b5AMK5MYJwXav7Zd/pGr
hQZ+yHpzRXMSxUyi7XUdNAZ1BGOgUphTosDav+zxSnGQ31SkRgBJJpEQN+h2KKUF
ClxCgZPnnBtATTsnYINU/XVQmMftoFOePbXVoh9YFAec89qXnamoivYx1WcYNb7/
WEd5zvf70LWNnooH7XRJmMmnMDlkwxjJEvrUINrg+ht8Z72OoU0Q/Dux+Byjgn9d
ssh4b4xVjZfgqWqLAP719ItyWHC3zegNCKi6Um1mbXwviGJcu0PEuz4L30l04yDI
I1B78EQFlT5veOG//Gdb5MDlH9IWowY9doE+0ncsOo/rYPsQWwpDDO0cXvXpteqZ
wlir1F1NQKSuF8MGbeSIw0fQgjsRa0nMrzZTSNESo2PuncERaDrn63Tdwv2jOg4m
f12KpC3Elf+DdySgne8MD266UkI4T2qf5HEQmEs37Q8JPVRNDfMM6B+2VpTDHKiD
oh+1el2X3amMRJF29p+5WKskpsHOSk4SNQpooNHIyBJrffkhTMCSm7TqVjJFaLv5
XF9t9sSdtlW6Ka4q05wa7LbdH08RUMNh7ffdtRu/BSmYFLiMtKEO1qb99rPaxw79
Lr+4wCneh85Qe1dI9seUvDAHHYlaYePGiacK1oIkWPecTm856ymCGX2M5eKlA1JJ
jeq1j0il3AqqMZWYB+e/LrRs3LJ4JIumgzCqogBWcjzZk7s/qDtT7oPGXCLzQ3Y1
BQ7UqcL2N5GVXLGUIIL5wzlHpWzZkwJRU82NLFKTRYCbKtX2nhPI6P4PPaxR9WbM
/hYPxG4LUncUiOI5iinHEEwGVftzYNNISk4LjWwh4j6vG/C2r2M4ntvpPjM/CauA
ExnpRpD1vD8Vq0XpxMBKoW0G/Hy/asJnUG0Rll8B4Pw4geIJHhdXUwhXw1DGJicu
oISOcsEe59gotA9wUh/wmoYs9GD6x64Iqi4lcw14uoqL3djVMkkn9ExRvBy0IbQ8
KG7ZuW46p+VygQWbHHOBIrBejmTfDOWnuUSPAANSC8H5+kcqrG/Vq6EhXrm1cU1t
HgeETwaelknYbzebxi6evLS81/WQBay3GD2EQWEdfTKuwp4QvA2IoaGpsq2Ndomq
g9VV2sSahAKexZzAqI/4JoX+WrZIkerat21kmBueojWZ3z3U2nq2ecqW00COlPWh
4PGcvmTC1wmrM7WlEWEi+h9hHbh53jg2hKhjbQ00bCrM0SG6PXzPutfriVcWsx/j
66qz2dPgiSP1TdxRGi1hBFIBjikFhPZBULodPv+6iYk2XqBZyUKWMVJGIVEuBV2g
s2eMUhwpyq11LFl6ClzliAwFvSvXS4PCD2bVDDUrsGyzGkhp8SwwFd8CxoabUo3i
3zkGOmjbMrptvQLfJC+ixkiBlWBtrtD/DAZMMWLmgsEaMwiXAOTudAOgM+Oa+ybz
EjGRdvcTHypStncf1ExEPV1p0/Pb/X7VNBEgjvVPcBBTNzvffrAzJDnUUfePhhYa
5sKzJgYA2DZlfjOgbSf2nwB0Ur2Tc92WoMmmSGSNTEUoRzGBH7XusTlYSVbvkKFy
CgVfoqRGU14FqQ4z4pFoomSTyVH26SO9DzFjmNOm8f62keCFhOJ+BkLrA52X8QZc
Mua9KinwTpESwSvocOJKTzAuTMfiLRS31hDumViE5CYRbgSleTAdIOAuakSS0m2M
yHMfPZs2LAy50vNHXMzOsTuh/SPrf+2xz+BqFectgqaFJaVj/2XAf2gq5jW97k0Z
y6E5BZDW3hoc6WG1gf8V5+q0Kfr6F4ljd9SqSgpTXfy0Kox2OQyp/asVX49kvfjt
YCwoWgZDF+IgV3zVAroVtaEuUDSajLXrn7gTXCiDaLM0Tcivj/sNn7UlNym5YB1S
qvUVhlQxuOKdn51c01mC7e07RqMDi/EVyerWXmbx53xEfy8ZHKyO4FycG5wYsMB7
xTmc4dHer9sCIglRpH+cDaO98lsLVE0HWe+Tujn8dRqZwOrAnMq74wDQY14r57MG
AgxpRZoTO7wxJ5sUMvLxHpix2RO1ricl4uhqRqVXAJ5gzlUMv2ADUfRzVRWvWsyo
aOYn69Ksk+LWO62dIQbRWLj4vH10ipBKAXp+T1PptYmbEDuZuDyTbomQmlSk97Yd
jyce2FGyNB1jU7eCsX3hmblbZT/dX2yDA2/YYuT7MaGsugz8J1QgXFGQ521ZM2cS
UkwpiIKjP2XdAh2mUMc7vAGeUjD2TDG/zkvJ+6iAWzFz1bCWkr9Juk+q8Hi+DkSN
RgtefOY2NKUyKpkZdsveW22s7rx0UMyAUmI6Zd6zMIc47fhwhJZhVdPbv46t8I6c
gVj5FXYNOhW8MkFSRt/Os7Q6AAo709UT4eBakJ+yXPXdMkFqOvabkp0S4g/wTlW4
UmkJg6Wkq1Fz4gwg0JhM5p7lD3SrufwOJ+jO8l8tzvkpB4Vr7YGS1FdverEC5thp
oXy77oTLZrBMSxsRu6lgRxkzWyCi32DlMbH98SoPGPdLln4dsLgbyRJzQoSOvz5u
b8gW5dIFTygzR6Tiqocxb0de+cde6uMhMXdBPDbbqotzYlcTnvFp6CK1KkvJtJ6Q
dDuDYs7cDvAHcZKz5Ljak5PfCVCr0pp3DdE0ItIM94QAtZaSdLu2yQ/EySIvkdOH
8uSSeyJOx/gHSPUrcwLzpNwcv7FgQvuqcqhfAnpKoP8N9jFBZ/rAMPUNwlpQH3OF
eM/NcEjd7HhL/CpbfiWyWh80JipwY0q3KrhHeQX+DDwEzKz2jWVIaf+QZI0tyfGE
Rppfjza0r3ytljoGAxzt0qFGQSOYU/arl9WVHK9yD6EWecmbvVJF9jjDwVM2tlqD
Fe2SwtqjwGAYP0DPjLayVNG3TkGxxwhAXfYNkKhBho/IdRkeLgw7dG7keeIiy7j/
HUStKrOxSeFMhZJwKr1zYOX9vKT6P5bWDxLRHlpWQHsC169X30S/eKmn+yh02de5
EQJUb5MsE3YSkEofUmnSzM8acfuE6eKlVFSbDadu0A40mGwi4vC6augvLvQqdgBT
Q1A8CTFEJFowsUXX1ePjV31qudtVHBH7S8s6fJHgnIf6SQnyHcr+hmCKL01EAED/
ieLX2Xdof3wt+c+A6fXFEBzofyS7aRHlE8AdSw845GAq5ABnoXHOafpMcI4TnXmh
TpyEmWYwiQ0siRBg2cjvdYQywqKaISIGnthC2/p9jI/A4M/mkAuokTPSLG8DIZnD
Ta4qtjKoaP0xpkmqjwgRsZF4iSlGlSUqrIN4fRyHjjq7mJ890KVcJmPeAvJmWVWE
ZmZAFAruu4pSTuW7m32IZrY/MyDAGAW1XeFgcMEab78OgRfOeiFYSiJ9d3Gg8gHe
c41ms68nGcmCF4BvWPJCbpkPjX10pxyDMx/Nysv7g8A4ntFru5jBnIJ3GxhiA0Gt
VyDVjdu25B7IIIVTSUZzj3whaaDUiNsGxkhovGJisSB9buy/RBDHKv3qB8QtiIoH
r7ioa6xgIajoGQmt3fEgRxcRzlUonN4Ujg+eMJ+ksBzteIiKh1rUOz5kuYxdaSh1
zlwsWGn5owjjWuBswopjEBWreEZtWpTxYy94wfUYj2S852Pzgw7dvmZFYPl20Gt1
HNSkIkP8LECStbcEcdg8pyw0SY53icewXBM6uZepHY6o1JcU7QNf1m4njbvKb52y
ATVJCRp/6iRLKDK33wWlRqzNsHkbR/Lk7n9DNZW7Rt4BCPL/9Ramf6Q5l9Foa5ZP
Gtx7ujCud0w3grlEuIyQGTudT/1Fr7/HQVVfVX+Rc54GR0LnqMJIRNTy/eedTG3W
oY7tILz9WCi3W25B5SR8tc3w/N9fTJa6xFjcTmBHmtyFFHacT/B8m2VMmklsqdTx
eaXVSElARbHvXIo2sAnN3PToGCylk6KuXQbjHPquINvBIMaNwPJB21RpHkxQkV29
x0keSLMEnfANOAAsNJzRSdUfH0bCHmhZLJgGZf67YjXD9eKlM3YHm7gY2MYkguEt
7BTC0j0VPfCATMcUu9+PWo3SsHv2IpnFGrsqN0kI/0knf/HdD6wMIP3kaqyvwUdZ
2Uw/du7QtwQjpxER9vQ5TpW14e+E1jh8T0jwQIOh1VtLcr6aNC3V2ZA70JAph+Pf
R2WmPSQp+skFIsB5kyIb5shSzR10M+C1uYrCt9L9Cg1fgqKi2YFhzbtB2Kyq9WLP
WFX9vmZMgdeiDZM+JYhl9fB+I/Qa0/0pAV8+U1HsOqpHTCY/3HZrQZgaICRpYMfY
/JBW7qKgAaVpJGkSarxlMTHC4+O9NUe1u4RZDm9KXtz7kShDAsWFQK8ZDMsKa1bS
I5DoTfUNweAd/MPr7sINuowXVHW20KPEDAHAT5CSLKS7bqHUAsdCmnTe4ekPdCqE
iZhqMgU4sQZy5TUVSNAizh7cfe9G3H+XA+e8w+U/eiRbTUvKgLrCgxxxYBpFjenP
Czp0qp2HMwmW6IaDBHjGYWnOl4eOOuVhUgzMGannTeuw4Hns8aRfsF+N4Wy5wXts
kE3RocJsBcaQr27k/CAK3ehXcG2NTODr5zVCy2nQvEVxxdzjbjMZR4b6FDnMuvq2
Ip7YWoDkS5yFwS3q9ZGxxai40m2hXKYbsvFF42xdLT6P0wYSS2gFWa8+5wqbVBuN
eEu/Dk813IMP7Vx9F9C1pXNWXaE9QPyO9uVvgo2a3vXkEjKBLHfAQLB4yhxU0EOE
ORSGUsrXHO/Bf+UTbkLm+fNpa2AyDzrHPCThL1OebzHWnQIM6o7vWCS/p13cg73w
VxzjmgNBjsmmyn+Ad4Cf646XE2XIb9w1KGkBHpyDZ0HLa1I5bFviE7A373+TB42D
2juj7e/TOfyIHZY1YwBZ7Wee3935LIBiqV5OTpYf2Au3ipwQlUMVkSbe9uTCLEg2
I9L7WhzbxwlxSVLDthgGXKTsH6erO9RbLJkezF0VVXZAQarRvjJpELmp9SvXNL7G
t7kt0Z/ktiC+/0QAXlew4XcAn5VflrkZjMN2/EmF6io6zyOXxC2QaT//HOCeJJwk
sPDtecWjRwN1BhEM6SoZ75eyYOC24nFvj2iSFX9nRUw8rC6U+IaPgxHG4gCNstWa
8mtpH9XQeRuT9f5t5ITypTBPZNyH4mlCUnvEPimWCIAjhbuPX15Ow4+w+SeZeKE+
AhfZyYfYZMn9/NMCG9WKW1yL7Lw8WK8fAOvVG+5Hvidz58cPbgG0c0omD9cnwyFN
6fHI73kyNhJAHWng6QQhjtnp4XkFGo7FXDOk0VfTBAOFVtMJdzvF1khu16aJYnG9
WoSdYIaqI17UiSJ2KY8cNyxMM6yBQB/edaTsjTvypE1szbGVjqNw/hTf2rfmphlj
frOEiCNsddMMehZSLDszTdAmF4jKbTG5D/1liRWDq5zp1GR6SStpian2BQW/OQ8o
xj/xPTdD6dARPNesY1gDnbuTSX1FQnd/GYhdCvODgdCMLr5x3ycG1Qf29ayuvuyL
LyBa3mlEzBpLhZDW1S/uiYhEtDUGKyxLMwAEZJ8+Kd4F5OJWJ+y0wgE0DLsRttnB
ieRff5URFjiYXtCUWRciD5TNKmnbaMLHCO9n4ENr/NCiy34Q2s7xiK+OHo3zjFig
FNP7FZ7+2gTQ+z6M9JnqJ9tlYZm4uTgLmqgyggMqUa+IWjiO6Ki5FmCO7zd9+rDX
8qQotPMxUOWemGnRW6lBGDwIC/1gC0UBvlsfziCsG2YH4dEw4VdTGohYSeYaFxhc
3aWQ3zoRpXnqdxijDsXRrBABSPwqBgcEfNcCFLpAcdu2ZyT27WYK4a8r1z8mgBFe
plsZQgEd/TErd0etwUOXnVbBJ7gOGe/oRcHKT9+tTUloeeHZ40OkK19l+u3NJH1t
u6udr9Mpew1bxIZUf05sBweaZJbG7gCcJ7NlRKWIMYUCMrXigF8p6gK3rU3kzUJq
RQGnMkLJCNmgwJkfZKPLOS0G/rT1vdaMY0jDIIQ40bRTdV+HE145tmlU7Lang0+2
T3U5LksIA5nVc4af3mQytQrUOrXo/UOxct+Z8TVp2LtmJEYpBndSac2Pn8zz55YN
srs3OhFZMZzUkCSHvB8jv8DrFY1oW1twzcUKirEgnKIZBWKUU1Sdu7VxEQvN9HUn
o6au9x1nCBH4FW78wyxcLZLXW1KHg+1vdJe0tMan6yKfw1c/XvbPSkI8w7WYu79C
UxOYZEO+aVLI5Duh+dAp58gHyyTUOA/m927nDbIYZDNNq/oxAwZ6wv8sbbTIBFTk
1WcdWPsN8VGepnFZm2IMpgrpS5jxsDmi2sM9tiBxyMB89dwKBr8SFsZusKP2gjPn
dHB7sBzanOh+ndeI9X3AZD7Hc/FOUaIGERcXHwuLv+miGnWB5MpeW3N+rdzwD1es
GJWCaxYUAvzTEaFzpBjyHCpzIg7/hzkmEzTtUDVqO+WTuCjjlzyhqnaAZabF5fLM
/+bWACnIb2p0cvzs7zvy5zL8tLZXnirRvqpPgpI+l4ivdMvHeiQnvMpeb5G5Fsi3
oLapPEwEmh40wwyK+SdTpmB6BvX56bQxm39O+X0DNFdB7Fe0k6TzCtv75DHX+OuR
pKfE/UeD72x901DA+CuNQPi7DVHjnDtysjzzIitNSg4DFLOeY1yUcG04ppaaX1SS
+93O7N6VSEA2MRR6ZNXVVDxKeAVtpMm7gg4MSFsKZhH24QwCINNsooa9M21ab+ra
vO/GW1zhOskXo0bj1IA+fa7GYsj+BV0p6Prl0vVGcj/DNhuBKdcshMWMi4pqLWwY
Qx/ANkNRExDCYAPhkNMaYkD0jUViso1f3okd3rTdfFk5alWW5V7HxIOW5hoi447g
0XAKje6VhqPSvOV+yZWy+qcU1fkKnOfo5onAsjrZMfzLS53BepYKQtBf01LIuKdC
1D9uNtyXfsm6lJOrNNSehBGW5eSFPvDJ8P6fL9zwwT71z9tQ/R/W6AkhdUJTC3O+
9bYoV82eQfZiwfC5q2lQEF5MO3vCW55NfS1kQprLAqXUa5zb/DxRHAhpd60lUGkM
s8/PgEY93QzOvtaCaD0wFK186MCjniBZ9cL538kCxdxiPifpHkPJ65XXepIErJT1
8yve8gdz5hjIq1Few1aXTd3PeNxrPuKJr3Evc/v3xShc2TiIQm2zybBKuTBFKUbD
/ijIgSXvjrgkZQ1esSX+6pegxQO8AfMZXNGm5ilbWVazy5IJbBr+iHhca27eBa+J
w3BtAWcWei41TJomGdFEcxixBF2pDOSc02BUvlLvCIo/AS9BOS/n9+V8z3yTT0iB
JS6bpax1lN7G7mhQUX/R0n84hxCsCHtY5cDeLX0e/aqm2z25jphlhvrYIHlJ9+6U
ampfoRTEXL2lw8Kdowc77EFlSqtcatU/JiBPr/pbfAyR+IW4hPtWUR7tof8jI41j
C0Lek1GjtTyX0IhBx/RyqmPioBpv7Tg1UGdiBNsFhqdYvOqmozUBUoPsLXCBiTTP
5Xfc9zVVe6fCfpG3WTwHkzUWNEhpZMfWo6eMw53SzQtgd+/xSVqmuyNYKF2bDpBS
rHP4XoMUfzG8PtREH90e2ELQekRRk8E72Zkf4jEnMSJfxVb6GyfoT7aZfq1Z2Mkl
rzQKDtAI6/vYk5wzxn7QACF2BBJLEK1hgT2oxKBS1K3yHoxxePdeu9ZELLV2t7MK
Q/ds3VaRfWnSkRNuD2GJJUXGWl5gUBeyQTN4NixP1qm8nFfJMuz5G6uHALfJYKb/
m7faw+wbt/43/o4VDm/3mOMoSR5zRIbHPf+AWIhCqTS2KZrTOuOJPlAZGsMQRC+C
kfO7Qp5Uf99bIN2iEiAQH0ef2MkriD8i2q326RT2FHzIkHsXpnZSlE4erxGCOftG
9SGfQH4VAglkJYC5lPen9bhrKb84d5qFppx8iFLFjs9q17q7W/kfYwRjvi5C0SuP
j1N4q42hcTFqdIO7irOwd2kH+pwpQRUwrwwLVAuNlpxMQsNoM14rsjV1lziu4djS
bxnCKczQS/3tt1sJQtBulfviEtcFAL7/adwfq0qvxO88OkLvJJzzzTsC3cVWjlnr
Ns2daP0LGDQ09hlu6d6Qw3BRy6jidl05nYuj+i5R3SUdA3cNXKlNVKXKDeskyhjJ
N5fUuLSMT8zFHuYSi5twXfz+DTeTcriMInYtMAMV7jSkCeojRr4eJDD4Ei2NyIBa
aZ5+2zFzZ/uJDwJaZub5LdYc2IcuoY/WJ+5XNGQq1E14LVHrkmbDkDobcIEBnURL
EFij7P7t1EY/Ab8ArbrKDSLr8M5h6jxQ8vbK/0SNC/4E1PoDHyEJtff8e0McJQbt
D0nhczVLvNDlJ9q9COxtENzRQdiFzQ0maagH8paBQuZLn4/rjlH2Cj6ltjKjTqRc
Z0hRRZJguvmbu1/aMb6Xcf6pnYVs5Ty9NlzRLIImm9PDMX3+yNfxzOnbjkYHEwhB
7WR40aC8VDuVRij3edFjKYRzAhkkE5KzMunCe2CROsQXwEe3V/73hcoLtikLIk1P
VcghAZ1TOFYVnEAa/AwRLou86LtfYyTveGx7ZpYVu6sIfCJYFeMICoRqjUHdPexz
GOvRfzqY3CIIdh7Sv0wUvoyyWledItvK1dpnYhveyN5f+wgATfCcZfDgcAHmS+zL
77oO1FVICjWeH1YiHjVQ4ljYpr+1dHiIjoiE835BGrgwMpRPczKKdd0r2YihLQ9X
XXzznn70hAE+Ud3cm2NrrF8+VAWL4GGuKCZizICtJNc69017xjkQVV+LEnc9LV2W
imMy0jVqNfKHxr3CeKK9YBVqbpvfAPF1Np9m9Z6R6pVans3vrKVHc3cYdQhwNcHV
701LCcn/hwBiYOHxlW0JP+lUuC/4xaeoorEWz3pvfmug23FQ2geFhqlOqJAipkAz
uESLl05TF3txbgjTJcYCQ67YriNNeizgwt4PjfBZMTp5qSoR5u9AMsITmGti3D/j
6BjmXR1EGTX7R/azyebKgrUte1yQruFG1YiT5YteJ8EL1JhvlkzRB7+cU1R6GmM/
FSdocwYYU9UFUakQt4fzlDZVpOzUQ4LDghYSUOamft/YFcOVAQoDU78L3m/qONym
3qvUm6LHeK2thpqBqkLqWPKvK8fM1ICPlNcKQRn+J/yyGIzgklYV2IXtf/EiuvfK
t9o8rAu34Gk6vfCDi3bvLyNdXO1PVQZonIit3AtFEgEYdoHuRg3HBgPTv1b0izAX
1M88UyoD6Jxxk5lJgTo/MuYBsynNvmWzwjOoEFNyfkctckgXclOTzkUjhQGFr9uL
J+lEmFJT0MSWbgYQU0/6lfUCcrJ5Gvod0g7OL7YURQtauijhxyID8JEb+dWUuhVK
0dAGueGxJvTWl/IhJ4KTXZip/M9HwRRfmW+C//FMo5oxLHwEs8kwhphpfoPUYQ9s
acjYnqzHYNhTU/LTGaagJT7xtccE9e4W5M1/ivk7qsRQlp0Viyf8jZkx0N15Bhjx
vwiQ8W+p2Qf6tZ8x3pHJLMIeauQYV9IJfjIF8Vh1KGwBlaXRCHSiTKdXEGzKOTT7
3dXKk65WGgD1E3JBRgiuTYX9fikptj7g/mPilMhMt4jPf19/6G9sB1c4lHjRjtCu
yKw5iDLTj7Wf5uTT5DXpVjKSWkgQEcmcLExRbkk6XspBEXO4IkGAzOMC4gvG5APl
LDwpD69ZIVZ0eOz5KLFlb1McisMT8LPyzxOO/09yrBMder63O4s1yPoMbjGXjtjN
f64k9/waJChuaP6oaokqHxJvUih0EwTw/pe9NqoLRBOLLEVuKvmsOy4bVizGmGIq
HBahMCy0wWK3l50KNzQnvKd1y4LJ8ZrKBRoxBXILLPPwK8NiTWV7jtPGBJl34Xyc
fLHvFvvuHSQ2oRo78PYXOBNdbVt+zRJEGHo3uhr8pbiVTG6Uzf7aW/OSsL/no0P/
Ev629q9CUPnGpB9fqH6MqwS3W9mup28oRzGY8FhaUN56DVrXaMyCuuJD7IHlgcXa
B2a5FkntQWQFImLwUJWa+HEAKk0H8yfwzse5+TEF7UOqtmn1OxF86qnGdl7TYd7c
V+4KeVc93Ma5m8TOuNkWm1oWknRMpNrmifWtiMLhPoEm6VPKtGhpy4qBh4yF6wpZ
/Es54fo7dyW1deCQRV0jkUmbYvis9T8wh9CdyX2GdNH32Am9BOqJ3F9U7blkzEiB
N+EohSwEV0r5HwbUzEM8DmPzy4Juzwr/zNEDPIMS3we5mCm3jYe9rzYvYYQxI2p6
0MgDLYJogVigpg3OzeKlBF3n2+LIniB1S4GUAzIzvwNOfrU50y3Kt0e3LavJPRJw
VhtYRAFoHBw1ieZY6qDVNTERVgXVQ1vkpBbSbGD+oYaStLNadQzJW+rvJIauh//N
SokwZ3/tHxTX19Ykv5ASQADEhcMVAO6MvDFaveCpLx4gvC4od1uphQ/gG2eCnxpW
uwK4F07j6eJTXbKO+4BqL4m0a2zl21Sujd/RgLjtG99eqZbgLV2Q5G/81QRfLnJq
DcMnlO2gbQBcJkPe5riQkgs2bRpiZHL4ckyaRO/y61H51QYkOxWxIqVaL0MIloH+
ASAW7OaUaaUpaPjntW3mU0qSfslkzC+q0KyeDPQbvHRbZUDMcOVna7RJrE3+ZAn0
ZkZ/FjDEYkkk1vSt1gJ7UfqyENouXVb63VjLs/iFfC79yiUF+6YSv4qrGrEiiwtW
uwFUOwX8UyEfv9D4kh12FHRZm5l9JU5nIpBtQIah/ZA0eVRqAJnSBGrXUzhGxmwP
/E2a9Vmp7B67ZANzZHfSYi5nkIbubDHyeag/DkGNcn4nPxdnkxrZ9QlXk1UjsSSO
tHrCek+5wbaIOHlj491NRr2YZ87prDFNcGW+Ide4jiz8+XjKZtU+yC6KJKwu8CTj
h2Cnmo6qJReSFd1q5F4rXUwXyig4zEPuwpmwFmGDAncuh0r9HCJFMp6pMD9osL2S
EUrugyFC6MWG1tWMcFtzo48qs0P8Y1pZzdwt917SSI8RqLcuUDhQ6PjN5Wi+VK0O
OrBkS0V4NZn+cf2ZOOsa/zO15rCTZLFmyPI08OTKfOnvHTeFYWVFKGnowyhgCqtI
PSo1rg/Vb9hZZgfzINC+VAnKLtjcl/YmOn3U51NG8Kb0uSY6JpDINN3b/0Y37Hkz
tzk+OHsgAzrge/dx8fMyvvov1UT68Cj+zg8N4xRM28C+5NIHsapoKiP9MBLCtf/+
e5AbDrI4ic7uGVr6JslDbSynqjxBanwMfdBtrvrDAtY5qK44m3m/NLA/RB3YZYk5
cimJNb22XYWGfI2Dmlq0JnNq7ilQ1P9bcpsHIidBs95HQTgFV4TlwgGl4IBBdJGV
O7QS8BmAwuGunhRnJUAHOd5zrHjJad9Qcxi7nfwoCznDtC8Lpy7Qi7lSJo8tqnNc
aFvqMaGAjBSJysyPZoNQbLLaGW1wLSTOVuj9w6DWgsXuo0zqDv9WACSM7Lnv1ZGX
3QagdphtYVDgNDj7YBtT9Z0850vkGtfe0vTn0C0OnAvvdrxs/mdcq3rAEfnKlj/E
al3bd3fah9WKE/FxARetp3RHdqn2oGVbhbgfd+Dp4x/YWUtm1dZ7pZ1+C/y6LTWS
4p384VnBAvIEjw3h2lCL9gm37WmAAVGFOqDNIIah6/Sw47i6Y+Nri654qLG5B6im
gALRWfDQdfvTzQs/VpzeJY7G3XTMIYq5lfflWwPh72SzV8YF+riI79g5jDTzNYuf
F2pf3XTChBc1lYbL8WSmMkiJohQpqT4Lnj9gM+1tc3xOC7L9j/epxvQuQpfnj3mp
aSlHI05oQkGEQ7wA+VAe+Ly9M7nOI4ya9FHSoqXdI2nLg9L0nKF4dXe9lAWlQRbm
ZGjzrD1qkhj5IVS+DVqBUYtB9DfFnqHD7Fm5diJlNXeFqtrLZCMQpnrkHcZkJ5PM
PRiHR0uVwvQI3AkKw9KYKUGT5uRDndP9kssur0VC2MG3UT3OsMGixO+7BJS0WAbj
NZpimoeBib37t5zjdPMX6KR87V1KKrRsus7fKFXnma9xs4Mt7WAfRpyGKaaIQdKv
+calgcDddKV8IIRfM8c9DF4MqJB2rU//1UqWCZUeEvlfRid7vso+aEk2lSNGgspW
Ukb08A2S2OccwqzTSPnabczfT6mrt0ArnfkJOb6b2zFoeNOdq+mhOFpXUkBbaMMB
gokgiPG38Zt6YMYAAdOStJ/oK0e4rlKCbaIBu5Yzg0FWW6tj87GC9MivM6241EZo
gbamkvt2T/V7SWPnR2BmlnMCq4xAAskoriYI0vpv9OIRxg/QoRQTMzcY9URd0eK2
JpoS9NPkN0A8LM7U3WNoWKWSz1wBxvjSXqH9mT308UzuhqWwnMuiqxo4sof77XsC
GUa7J4TREH4dmzid6dnAiG1au+py5K5GH5fPLe3cOfA7RM19rPxlWnuQ32GbnuZx
+IgHCMr0FmbxWh3lhjfAIcXS1Pr436DwQgVBfIewCBu4D05vmbtI+C7ehqgrM3Nc
weqb78Rq6nJSiSFhdem+SNhWeVJzPPzVRbzW35qCctBZiQkrgoOBGTYSlgmyUNWY
lFQdHRQHa7WVqMAg8vBACPO0+JamJt3XrNAnKc0uzRVkMpnKBbxT4SC/XrUvXcj5
e762yEw3S9AwvBThy51MWZyDrGYtxwMSYo47p+BLXQi0RnsDEKGAUI0D/Cy5wM6O
Yu2eEKprvpLntk8UURhb6BCJ6mjwupIfS+h4UEL9R1DZMuahevPZfwceRG6oZH8w
Tj8tR64n202yWKRrZElqsQ83XYDWbTNC+HJ+bxVh4BJVLqEfdcAsFNDw8hhAgvA9
9bDzMzhF1z5kal7nY62EX4G+4ffwil0/qbv4Hqv/GF8E9mOK/upozQqydkxw6iGx
4ELL68n59jVCpFeycQrwPoMHESRiGMlyM0PgCckBTIXr7B6W6d5keHHAcQJXNBnL
mBrgYMMNB6COB8sSJR73vJHSc4jRt8RxrF+RUZsIQDcKGHaNyvPgus0782vFQjbJ
Qx/Q/LKCGoKbzyUBZc4YT70X2k6hK8z1xs5DSqGxGjVAkN4oqUO5xQjb86movmAx
v6Z+5gaUkP7ZQCSd9GjmsC8lY7rW4b6CkMYmygu7EplfzBHouViCfeAV5VSJAkUP
i62fDMwSmeTiH6jTtzRo0uGpchphUjBCVeR1THfsR5ozcAJc39uDWApexs0MbcRO
BaBcHMjJZItEJ7CzEqSKYez8lQaW1Ip+bKvtBkjdFGQ/PHGZ4LYucUoVcFRx9AeL
f9+ioiBYFtNrQGDr/+D4YMbaF8PQTeGiZFpHMO5E/tzVt96w3WrAxaMtNlCeMwbW
dglel9I50EEN2NlRB7kzlNLRUmupvYmObtXa5hrqprUPKOO62B493p1SWaJgdqYF
OTOWh3qPrP6aNKroOCP1/YNNdNS8HyUjjqwZ2ntqfQ35mv0ZL0MIVsPGch6FUo7P
4seSH6P4U+vPAGPIKmrjaQFl8AKwCe5G6OiMUV9LjSlcgN6v++HiVEHihBdxONti
s64NntYtr3neUCSVF23pmvF6DIR9bjWt3n9x/cnKek+UlQiat630ohd6XE4Tfhef
bkrHuyKmoJ6/ORPp5iYizw64EL0UYGDABuiZogtf+cFA4YeRcUKcq3soItV1ZZlO
MFgnaIaZtifNIntzVv3JkTMkXj57TU3y/dniWxEPnkv296xB4ym58belfT0VqmkM
O6hYY+pwvUYbpZCEa262Z1iyJ9fGEsy5hLW8gy0EOnStUiTsgIDz9cU0TuGRIpih
/ZfO8NzPVBWy/PxHo6kXAaV7+jx3FmeO7MVJXolmobTeJ7v22OQ69ZRMq1P7yGxX
jNhaTP8r4wwNRBiF+HYx6wZD1jOdNUNfisnGkYMIcZSArHvJDOeaQ4JJtANupxll
Vqq0uLyk38yQYJ1Tug6cStg/K8kVvOAm5jGpawjfPNCFSbs+8Z0+MrV9QkuMUEoT
B5ZealxM0ar3hItSXOaumWrN2JArGv5cAf5fyoaZnMaCTpjteFA16CIH5WPOS8kd
lB0A3QgmbN893+LbBgVJ7n5MH1ZZ0rW7+OHIBq0tjv2vl/IIHnLjAgGUYCwLJw80
BAONZxWvh7//JvyaRYCV3YaH2vfrdL/Bwzf1Gq9wyQkJlgUS/+xrswp5TPbQ7HU5
Qo/fX5oiMU/AmKFUqj+x9nDiUE+Ty1tR29raSeLI8ycqgb+WIYz8tH4mSCafLmpH
hNi7egsTEbKDQMrWvLgf/Pe9FAAGxACgdFRF4VswnfbarihW+FLx7s0YBjeXOCQv
u44H1izeOfO/bDFMUvncPqDEf2P8rOfXYIfCyT+OIh8awNmx+7+fkKhEdB7roEiN
Y51lcWb+773CeJgaJCzGwjigeUO9WGbrrRGrfj0rAQ08uRjGSUDF3pYYtczvtWa9
ZAYSxEfQcjmG1Gp0E3iU8RcOKx00fyTYrSrWPEK8wOyOavKz5ZgW53EJZQjgCXem
wzc/X02Ayr3kCUsIDvZW+/xJPG1o8aGxQZLUhHhPKJC5nQuxvs5RIjgN+iGkib+X
UuWMwgvhtKu8l7BWG03ev3WGM4zlJ9FHNr6gF6ZQeclkXdKuYqXOTcIGzJ98YuB4
ptrpwXEPX+qyIrZTtWiPOCQOisfeske4vtR0iL+UrKBPIzi3hJ77k+XmBM9ZXGgM
buusCfZFNLLuOew0ICKu669hzPKeBNpRM/YrWKmA5Pks7w9KhCPyTr8jR429t85o
R+5rZUIWjga2G53KZAYQgb5Dnw8Xmh+3HwAfKesicQuRjiTh5MQBmj722rKgPcaD
DGXSi79L5PDzc3+L78k2bN6qUEI6/5kq8Wkw0Zx2Qa0MKEHuDxMEeMfnYCuc8j1+
hIafrkUc/5j3y2P5X2gwO/VSoR8cAhc6BI85XIU8ltwHcDWucrhheGTNzOkzaW8q
LMLPLP+EfkeC1Ts2YTiyt4oVRQiHvAgI6VHfQf+QzLXsT98FL25BRC3Itx77wXTr
KLWq1fZcgIlG4hZ7jrn8ALtYOlWs948myMoJxi79B3s5gHfjx8bev2OGkVLQHOJA
1qcH81iyldbJE2+Luwzlq+Qcj5O0BPFIExkOLAVrKMv0RYSQ3TurCoRe5syK/2ng
dkypNBh/NCHQosIthQ/M4yzqVBy+PLfeRhBAPNBJAVAsqHS5Z0FY/XJ+mFbDc6HA
6e/pQnNNoQDMy6r7i9kwTQJNSdd+tkxA2xS1J0olt0rljVTlSFpxPgD5uQS4UxjF
ElkVTVv3Ce+Klo++gdOQKglHok8EEnkHHOm0rrR88El1NB8Go7esGYGSjesln1bC
qku8TWRRR1h9ukB2TqxAklmY6rGWwdrfPyeTCNRVD2Owpt2Hr8rHrP8Mo04JC/fh
zFivBkmkR/yu9o9P/AHS10XcBK5LvkmV6tTg2I4ore+/LLXIBZ8glK9ezBDsU302
e/ldTASIVazug3+XsuggGM6zkMeE9iNcOo/yaf5EQk/nPSnPx1f75n9YGRS3w2Tm
2Zw/hSdfQylSDvTq4PM4waKhmLMOQ7NTblvMhnRfQy1iYDiWjUr/eZ9w7Y3nYCYW
NnCfQHNt1WEu6/lJAqsX6x2R1hiJWaFTr04EQwVDRU2YcP/B1jMyGPOA2YJIxnXD
HPxX32Bu85Fy9phcqGE1Kp7UORTrDtupEu1Rmu3a8/4O/p76cIL0+e2qMjvfLrLe
duj5MPF10Hr6RWikByD8ob950gliYAiVqnsOCqpL7m6m/c5hqFhu9rLwStKXdYm/
4ejpgUcEPlxDF8IuYdE846jtXGWq0pbXtFXRqqm3gmnXBjRBhnwURTnlBPzWQ8vv
q9YQMGdTmRFRWrLlDg21ibOKMz0RyGXTDOcYpZlF8+p7nkx6vPyK1GNZ9rAQD5+H
wqAVn2YRHFg7kYKxi/IZuqcuEflRPmiN4KVH6jw9pJPvEFJGjkgRUZsTzQxYNtvg
+iozjfnipLsUUWnKVdPQXUDsKcUI2rtXeOLWmcQz/JteH21OL84djPNeRc1IyitX
XJ9mBejwEFgflcDBZn4CmUHkJU8VRSCYAGd40h6vWKuHr+m6mswJhvxvrKdRoWsL
ZOmopbzw6OELH78wtW2YfIFd2J4JnqutPqmeeeJD7zd8Ekrvmbew/XsUYb9a+C21
jmu8ETZwknXi4vaCyxF+jDO77WafEx/4R+EOwPFANuhaT7u1RZdjNSCzEs6P8mC0
aQN9BNwlNMWqZm9J4Ghw6gPkREqpPqStBOrjrdnrTODq9WKyIKkE/sr3XBy45kEc
apsx/tNR74Q0ler/cLBUew50J/chzC422t6dGpNxKtbRwI0R81US0CCqG6CPHnCU
r2w93RQiDi+UKTkE0IHMMdbs6kA1SZArwvl1JJp71tAxkDUwerH6O+3AwWoh69Rz
qKEsbqzCo089QfqvP6DLzRqeAlI7V1SvKZYaj0dlnhy8mxJ9UpP09bqEX9Mp/wbx
rLrP/j3aN2ICXDa0HFnN1DAStyryrKMYkMs2glsbocyf8bdCxVPWhXZnSr+CMwwD
kKBkXaOq0vZmiVsL2LUMZIMVHZXVOuSTLVPa/qJbq+Z+XZWs1xiNg6va2kN3LrCD
CBoR/0XRbbjVT2O03ghdlJkW7Hk3K5s7dImKsj9CfAD1yV8xUS340gzkBvrllypS
oOOdjDIONhF/9OKQEUt0Zge8+PtU0QtJ10oeyu1aliS7Zx5V9M8P6Jr2TLZ9a7JI
8zwzey3t4ZZj3v0IF17zy+ng74Gspc9VDL3X4IRf/Iiv+S8ifBTfiNUnMFD9B6OB
xWeapmhC+fWWCpzlVWfdNrOgayDNGmHjGVSFbTE0bWcF01ZCO/tSnnGqacmLhY8I
eCOfrEcUnXXJVNYBtMXSRFOuN/Pufhss8aN3Cu9dNpr5Od5gdbhTRnsv6vOPfDmj
S2c8slheDSZHPpo37DhPtUYau7rdAh8Ib1otC7vOgmtv98zdA/6RGhFR64hLjJln
1ssBD2j4nNAxmrkxeZJ00Hvw/d16O9XZd57iylf+VpOHNCFee3HkiaHyZ7y2S+Ya
eXSHbdL1BzP3GMRy1s4/7rXQJoPoqsG3UbY30VA5dfXqSNPm4gB6qZDYBjbc106b
HRC7vcBD0AWzySZs4rq9GOixOzzST9dVf6X9gsZRk4EIQvwJKx6lxcz0wYOvGhOI
GNaU3MO/CVgBzxfpeyx+eyM/xZgnl9dsUtPCkJtKTP5LeQMoKNXy03RISqjbscd5
6Xv8AzNY1Jc6K48CK+O+eOK8HgHq/G6ZQTLBzpsQHtZg3UpNgw8/uOxYNQwf06Yb
AlAgkGnO0awk1+cDRz/x6OOfSIihkFjrkPTFXmdtCVl6W2PS2YVkt2knDfni6fBr
TOYSus5bACxqC4U1FNAgmzNcDMgGqlDD8n2z5v98W5OA5+vKtjr9HhrR+vygHLir
ysDgpNsYfXYNcp5xfCtDdJBhC4wOOMK4WLRBSC+mxuqeXifJJ+QBkRrvBJTtjpij
J7VIrvnV/glmDHeZblKvD6pPRjy7i7dkCR7O1K8Vvcjn2eqycA0qqNox43qBWVCA
vValS5+nr3E4dbJNd/7RoFqbuQa8oaqzNuSqiibZWJEBx1JAjz1ZOuMigzn6RVow
iKC+GBJ5Jkk/Onxu//BGJx5W3hoFRtEZrm8I4/nGAU4paoKaHehqze2KLiJgQNJ5
zWIZLn9M4QzV114WsgYlBhpPZ+JhRXwqX5jNcJrRO0AqcytU6xQT++5g5FsuKlWA
dVBEc0gd6PsDSYtF/5iORcVW/bfJMiUDJ/OJAGB0auah+ReptDY4T520vA727FYL
b6eOEqGRKGnBspeRT4KY0Eb0Mn4uExgzasug66wHPihJNtyt6jlVEPQ0wP1DN2gd
X9zWR+9o9f0+tKAstcpj7rR6qbd+xoEbbzYRZTkM5PpfrmRjEz8Dy97BMBccqR6b
0g0c09RMfAf8CqGobMrFZYl54+0qJRimQsbLsgGMYkACsP+AHX7ahNhG1SgNa8YF
gNt+7nSdvMizXg4DDgZyXRuXEsq857Doh0CJLvFRyQQKS8vh7SpzSuEKeLaCPSO2
yp9UMHYG9tzaqPj3M2e+QujxlzOX/eub0b++tNE2wv5EqLbMzVN98DV1GCrzvCoa
lpmAkJCqt26ZLbQpPcmAAeC8U6jQFjEOmLO7qj9SENkX9h+LtQcA2tNvrGznQ34N
8XUh0vxJ/ms/f4FbxfjHexAA8yvEkTgE80MRNpLI5yHu5KUaH0TCX0zWEL3UlkMi
58/4g+BSmOqM4iJ9PYu3jKHoAGyGFUTEBDYn4KA6vDmY2F51Pu9XOMDS7h1tERsd
2cGdmKypgHl+CFOXl4v1KJkQzhrp44FLfGdQTsnpRYOBRAZ/IGPGqhttjL7Nmcp/
/Efv7/d5ZTd4TgSHsvXmfqS+vH8TJqGskBmQog5sF7HZQuB0leEYNfPqqIOdsK49
zD8Gcq2aFE71pVkj9MT8mMaCUNfsQnLHS9xSGQV94HcomIo99HtdOirHOVoOk2K+
mCMrCyoOG1gqQyGgPn2klkcxct584/wEUkp2K4z5gvqrpk5r9oo9KvSqwzBkJU94
nyxBQdaGir5MlxCpSXkpWk9GWjwEJn1EX+FjsEpd0XOukZBwRpr4AxcDVRHZRRcC
znOin+ZtjF+rKYrykEigXoczhEkR4EXpfSgY/YjkmPoiCeQ11vEgHRgMf1HEFmn/
9Mha9iKpwuqoJcaPIh7SvuDTL1hcONahav+l71vRwNMM6imBF4pC0XTHOTq7HvT0
a8dMd0v+6qjBXDCYvnG9N9UMsPF/UL4PqLuNbEtvjDMDZwvio/puU6v8tETZgDhW
nmrXEx9jgrkAvxDIpcuNZpm1fXoSI6gEYWNLaleirs9J528DcgcQAOesAZklqFRj
yxFK5sukx+xHeCRi8A+T801YQkTF1Ix47Pc3knccCW4iNudHoBzrhquUt2TWxA5/
T17YLY1rcOOJA0jLInhNBTx/jaAPsSmDialMl/5ovVWn/r1eY4cXk7KQemPMNI3d
xJcfNxRjWBs6Z0Biw8z5wD5n6Okdt4uHeN5k8H74CSr5p+uOGTcwkY2ZDdypn1oo
yj969GQN79/HeBzQNEBohs9fpNrbOlz9eE5r2KE6TJi9iAnTtGtFiBYfwvoXiA8V
EsnEV0WHXvkg+Z5YsC2S7T6Fby5VzniBHDXeuSGOZUCUz0/scp7IF9k7jYpbyeEd
FGxa6byDpWbNa5Jq3JfCMcMJgoevMIr8V34JzJfcOF+u3SeoOI/47By6krV9MkWn
nWn92Vx2QAfRDYKr96K2KpIz5BoHOITidzjms4+sn/ubQ7866hJsDZpnUJF0YeQD
fw31t0F/etlTGAmkHaFtsCcKs9VTdkB5nyoHg5CCOEswL/EpfyFhBfMMmrVJ7ss9
GgtmPqLGBL3VA2Ttcm4pCxKMnj0ohnZjFgDMV6Q261FxxRGBGBDfTiX8lWoJVfCv
50W1VjmR4PqYMAdMCAL4jADbhaWze/rPaOrdJu1Q+yxRKZS8KNWIx8Q2G9I6kiel
k8p/tdB2UrtDI4X3RbB6iB1lPYeFTSlWUk9ytKIuj4IxxXoTKZzwSuIt5nJlj8vq
fup6mbbdyIFpuwnCmrBSbNG0bFDCNh10r6bMxb4sKq1hzRhXaBXGdo0eM8HusCMf
DLau1KeQ6ND8L/u18jZQnJMShDWkW/e0E0UgwsUb8j2yicO6TE04j486aUqWPTiy
NqZrnmCINCVwTvBl5lOXHgTsn7DhgbKlhAtUpLyuMf9MYqwvNEEAACyIK98ZZYJG
mhQUM2ohqtSeClVqCII8cP/kP8S3WJsiY0SWSXVhKX6IewjlHQRUFZNwP31zPyv9
EBXRlVwF2ZA4RV0ULyCiosCVReqO2LDYbIf0Yt6EjhKi/CqYX1MYyD9KkvZJglm9
GlyyR2cz7ZBREciM7/iQ6N8gRFLb7IrbLGfjFnztClxsurhksWwTHg+lG3cs9rvb
fAKmegv0eXdgWD/55QjYK6CMYePpYpFRuDGmmWm8AUxZhcNndqER+m9G+Q7jlafj
+OKg2AEyUPCdDON2bAOHjebWJt3iR771O85rJwkoMCPz5fMKLNeC7csI/rjsmK48
TTGlzDfiM/tWjqgc8tZuNlGIosxibr55toG6eyyI9rkTZifgVOYDG4ucKms5E64y
PmoMtWDtTe7D8GGtFMU8G664Nhs5N+89UuKeUD68Flt3jIBqv3vDdWhBckNib/pt
+jD9xiG7NCW7avHeXteGfCNc76VA17Oz9mZWirCF3oVlraLpgfCkHQCrbs01tJeE
Ax1v6PaGXz0waifhwiuMRyRrg6Cl40qjT2AYIphBgLg/O4kJ+oyu+etk1h7EF9bI
WVKwjPP0aCmrqFZu7jXVhpFFdKEH4q1iOThtsls+85ao0232S029MibevbdXqHzO
XyQZr39OZoVue+HfIABAx2HCg+JbRUfTBg6lJQZwmougeF5+Y9JN/EEQb7Y96Aya
+Ooes+vrF2kv6cuEuPCTUOizM8962ThT059SHdNBMT6/MImVBYxyi6H/u0B/AUnl
Qjp17GbkXZybbLy0cJY1X17eUgkQ5+KW7D70hRbk0nGum11cg829dq/AMUlyyXyV
YVaiTYwxL0rezddSaC1Uh1cN9hXMg1nd+6gWYVVhvg4Gzik6HFsd1pbDCWYKhJp2
XWmeUEbYVe++TzNTVzVg6lwdC1t1YsDHz0GJY0GzDHH4vMo2p3PEnmC16ktBpfOy
ebn8fOba+NXome7hVReRRxgniuBlPMRk8RVrG/Y0QSvannwjp3w+tPdpI/zUv1kD
8N09FRCMxr7K2siScOoMzKNRa+37SoB99MlzqKu38Ld2sPtYBADcHcQC2m+4LtAX
6dmEN8bq2X3+4Gzkrogj71bw92oFwPuWaSn/wle01i/w0mGXG21cDt572DRYytvG
Yx/JHPVj/TVxvHYWPMlbEL+U6RxsZLOa5creKyn6qauwVKkmkJ3k1coh3N0ETPtV
DURIIS4/pHM6cu/wElokGGG1zMk40ZSKMA75OnV11T8x9/afqZ5juQHI0LireHSt
Obi8C2RSbHYZDUlY7r6BnA5lU/F/n5JYOc4pGwtnUq+pSmaA7mAXEYo46qStL8LH
J7gWZYsRwjK6wnqcWK3lLJoSk9dFXuvc0nN9PPFxWg3s02icL0IeflskmhzcljuF
jTjfaYRk9PRyHSnEwU6yLUzPKdEP3gFHIk/0T6o37WS1D+jSRA0RnUbxBv6/0lUP
bk+6FfpBJma7gqlrCHxF5zvkY3TzNduw1AuhPWrVV3x9Y7F9akMvSH5F8v4Q3Tle
uLgKGeIFdw2GIYg6a/OwacIa745BsFZ30S7BQ8ILTsvY9wUTHGyCKwyOnQiuW62Z
SiJjGIFj9Jx+zLUy4RErHSExeFxB0DwJsXPC2na0tuk3ioXv3PVjPBZIuxqE9bAp
wh5efqcNz6sfV+oDpnJQzJTVmK95LluAk7UtNaCradefjoQ5P0h3uJapBSuPOPJv
8YY51LVQuCnuKHfLd3sEpx8EcJaYFt7F7VzG65TRXYu5YYXumvpaX06TFWXy71sy
LVK5XTvBWpaJcf02n+PU73+L9ywL0bcHT5tyP6kBemHvhxp+NDLR/Wlr4NIorchr
ArIGD4jn2ZQ3JlROEp/FBhcATqaJEnsN9Kp9pPgWnVc2RIn2AaecVBHleyC/c7mZ
KlHGYsEnofjFIiPfURUlEl2BuM0pq9tpE5RbJWsbMOHR2vAWqVWZUysXaUXTGil+
yLt79949j/w5anjMc+3839ku4AuXEUK/EqVVl0bqK5tlG3ShCE20t8NZ5DRv4Ndq
YuucAP3DAsxLs+qCk1eCAYXHGp6dvS/DhAnHxblmQueFL069BT186G6zlNz/h9ty
IdhnR9m/xlBNzsj8vMyluovz/NUWGRZ9ELC4RK5Skhtx7o9N36Relx9wjdni/s5I
NYXk0ZOiXOEXv13fkvhil8PkyKuwmLpEHHdOkweHFRXi8dO+THUjLoxjeZBj7pn8
kkMsQlQLdAFTBRs3OGBc1gwP9Jl6RblnvrRCMVaYS9exPoJQ8N65sk3KABDUdOOG
y2piul4vgEggtt0a8vN4iRGIoVM7nWV/ERrPhgS8zXYQVnCnzTfpbYk492hDDKB+
3ZoXZCa6B4D7ooNTZH6WbtTjzGWdt8XwFN0Dt7gVLPnKd8FTGI7fvBVGeEPf4jrm
8hC0kIa8Oi8mRJdN9RxkBXDjTTmRlkqZDSW/k8X9sjNad1AzhEipGEj/T2DduENj
keztWz16mDgJ+rZvQNQkFg6Cwe9awOTA5UPBNedLpQVvwDmNielQrDS63RVJ0XDG
1NMPjAauOqkolnkMmUQDedAdh5ZUEsAObyfdYliw86zqPQ4ef+jcvPvI37eqOCHq
39b1jS9WYFRRSNH187/zoTGD8LY1/X1e3aJk2A6f0pYSwfi94DQIhOE33GPXCTAv
AFfNw0Inu8QOWxfMqeNZD9F65lIhNO7/cGVeUFNgoZDcyHrrrngHivO3W3HjDVaP
oaFH/FTMp+8PPHINbZBl42j+HLNKVMO1c+F53oJfYLePgebK4t5gNxn7erWQIXoi
EemoFflnugPgFMJBQPT1nWtXD3teIGhttO/tgwEY8VRk+ByQxiFSddhaPob3NufN
d28pBttvY8OI60NxFm4DoiIsZjpQgSb6D8P9XLu8TtBVK3UesERizttqKxNvF43O
+Uw4/h027TWcU9DGqIPW4jL75SJbMdy7sK3uHF4cYgT3Eo8PuuN5fevLkxEMJ4V/
8ov80z3LULjnBkTwOGaoc1nRjuZo6jAkDjdozz3jnQyP+3d5b6czWzpKOm0/zWDI
82QnGVFrZaggzY8TWIk+47fU0FnhiKTSRjbBfO6WD0NXD9xDDOEi4Ja14Pb/ZRZP
jQh435RyCJJX9fx5yQQVkuhmGy6nWRFjgB4n91CM6vRERYvFkuLrp46MizaeQL3L
qhUyMdnMBnji5QmORxarQIV+kcA7AvS5axaU1XdfC0ttUYdl2qNYHBzUCGpkW4CM
A35bngDT3g/5VuapdWZhHtYHDEdv3EFovgaw07wkishdqvd5dvvrBeBl77aF6YKe
jhUprz8+LtOhhzLEm6j5iZoX0+zDcPuI0H/Wn/8CyjDCzDy9NTsIJBiFLqFnbenm
xs12s3ztXc7VKm9OjfO7IGtCFFLpCMy171ucLDwDpYM1rPWYnF3ngdNov6iVq9Qi
fPB5ipzrqWwzdsCMuVwoSZtBMe7lE364yKxhNn8+GOerMqvJ6Q9YlB2QX739UYA1
c1tXVmdKVqj/21D3myE1aQ9oX290h3DY1mMmPLpJSWwqi4hZSlzj2MZn0Pyccf/N
3nF8mAXyVbH4jWt44ramOgof9rGuX0EdhfnQhzQxoVKERMllNVX80Aou0t6SJzz0
RVsAxcYf5cyfvsVQ+cNeXXD6tizVsfHg5wJtZnpLzl9v0iESoCVJzlgm3SACrAIe
61ul1i+AIC5a2wMSi5QOwbTI00RVrVuFGcOaaCoAxdVqLKZp0g6A4ef5bTNtkK7g
1yMhcNxz6xLijtPF3lbQKbT1WRrCunXUNvD2gXCj4uo723VkV+DwPFTr9oq16xl/
Pdj8fTa0pQpuRO6qp4qclIleDGwd1c4pybxHa2TK0MISVjn7J2xg8+TBmUoag7mR
kj84/g01naA8EvHGzq8Ome86NQnUUf2DF0dJl+yH1YYQJAByYPVqTidnrK8nOPJ4
xZDmvTLTo9mIqqwUnj8iFzVlvhnlWZtAEnG9igasozVpvKgDNuo5bbK9sYJaRrrP
smNcjqFzCZhUcbNiGquEgMXWjgxwbRG9qfxSLDB6SAy5bYN4WiJ/Crt6zGT1z3rc
YdHfwxYyBviWsnds4vPgASOnTk+SpksgT/kfJVRjKfDUm/fWc9v8SPBNpYBJawh4
7JGWSvbHRX0YWDEuM7tZDurrh5ILlSTLzK6N3wanDmz/RAmJ1o9/7hOFQhZh7EL0
NgUULZrkdrFkTDMV+s+1CqqJ9507PCI753cqvRkxmPO3kLpD7tpF56PNC4jhZ/4v
rwsfrUNqVx55o1jMxyh6H2XjbY7ysH1L7Y/oVVGiaNV+Li9+lLepYxXBzXBvXRkL
KZ9xY0bb5pxEAx0XrZt9avx87jKFTU6+r4X70J6hKxXMJ3AOG7xcxN99dlzSvvDp
IeqqyzyUSxdjzy3lMOs5rhV++lKwFTj/h0covqLNovHx13q84UNj9HIXdqsyVZm0
LE999HVfkHs9KOSeqtM4MxvxTFBYLxez0bH3QQd0B7bWcBwL+bJHrIlccjByjpT/
UAtjpAMjXyXgT/LMXUTlyONvbLiklk6LwHKQ3z/ySWb5S+jVxD/bqiC0gbyniMAc
pc+tqdc8rb9Q8c9iAAXe5iwTPkZbdV2a7345GM9JBWeNo1gkUBN6BHTm2fzoNvRl
cU0AXb6OGWoGvcuRdYVvqoWq8gzyINKrz4zMpY/O0dGkrJO4Z/DNtSpxqDi56zbk
yVWsOVxIw/ylsgU9ka5eh+ncp1bBT+QKqb0urHyeNU/TTxgOivl6LkelxyouIZlF
3SsxivvDlbvcDW8al6ucBxRUx6rGAYPTMNOEOt0wppTbFTfSKrjZNrptJsXFrqok
/wj4X+COk+X+W6qxmNuffqx3uXbsjEClPl1CK0yCBNoBBLxLJgM+Pr0lWIPNcM/S
Kan8h236kO9iWGDEzZiMFr9c/3CvT1YjfpwYXBMJ1DG3ouRIZMlJeWnNo/348Ko5
sVBi2msJbItOSI2UE7YvQW2YA1JxDzFLJBNi2UWNjUdPB9SMRcDYZg+d6C1oD9ZL
FsL4y4W/orBdcnJkNuTBBpnZwdqOxfOulkSEXIAX8nlcG3g20WN+4U4Hxs/a0eKG
oEKWttoJWbEPEWDCppLRZuIoEkiNhP7b6GXpZUEgCeKsWbPsTsnXuhwEgbaxm2Lw
oRKfNAuQ+utVLrbfBEpIRvWyATQj+Gk+PJGjVBOKte9TiV2mhKIxkZRJB6SCVhUa
jyLXohWizcW8cOKwilPHPRiCNCyOjMZWIVKRN69WzhKAMEjZhVgT5yzEEuaGmkkO
uVYMcZHdlB1QngMI7hXUhWltwwdrcTN9tdQ7JxPBMABtXgNpA8By8MNG8zr0uNJK
5qQaT2yTCnWfqtb4KHU7JFfZW1lRpSlTsEq2CXNwoTPfHB4AHpJvZYSGO+NOynbu
basnzwYm6tksJV7pL5YooLGBqVn1rOYj69G/LarTfdPe1qIzgt7CEKr8p0pHM9MZ
DO/gidFjwUM38tC5uhGJFk2vX9IzyOJb/2RubaY3CVlxahZJakdLNyBB3p7/BET3
FZuGPd3EI4B/GvZdXOfqyRpS+yssoZeAy+/eE17JnAjJKnABemOS1FGpmjuj3kzf
EFZlEg0LncOx3f86FGFySg1yM57i2IVPXfl91Rv8h1J8ZPFRYLWzeYNqvl2IC+zd
MLwuHlBdYYwLLFa4W+fZIjePMwb5Rq54buP9I5XtiYxX3Hcz1jOkla30XIGrwtNs
s17TPwYFrZE49vJg5Dv4Mb/2dkwszPRD8PNsTDVyJ7bcokCIh46pkG+u2D3yV0LN
m0c+BDmxaDKguLa3yG7Ry1ZjH2TYyjm5Uaik7IBGh7iK8os969AIYPWNhi/0wm86
nY3BbJQmyHKih/JI2irLrtXB153vTPbe6K+zU0Qnrm30sD5uWN8fMipsjC6nMCCY
h9b01LEuDJBX6UX75mfZJGtR0NBeBMB/hHT+4ezK2Kr9bdPQSxm0QSrhIPZEZF2p
zwVuLBcFnWW4M4qcLKbqmJ1S/JDZ2TGGxbo2AujPOHXyu8qpUQAE6kIjxjNEiYBk
Uk1sOKW2fatioKLjpTW7Vtt8xYRH06RlMYePhyGxzeQxhKjG2lVIaEXdBapybjKE
e4ayePG68dQcJfq8ihp1nnLfqAbl5+uOUdrtuMX2F5WSLIfUxOiZ8mKowZ0xcqps
iUZCtFGiJTAmrzdIc3KpB+g8sID/vMHqEJiGRMEPHy4GqnPhevBnMOi4pLROy8uG
Ia31053fYHGkyxozp+GBw82PE6EyQxnoHrt2P6MO6Br4XYjRKIBJ24rDN09KAiMB
ShfuZKHtvuLAL8Yqs4znHjR6V9+e69xUPH63QfEFovA87eUscbZ3nrC1k+enJ2UT
58JtdvCDhPTamWulMJ0Pz5B1l3rR1no0hleK2D6B3owAcjwpA1z2J7DNlWdMMghy
fDxeH48Mzw3XxvALeHgfftNBRSdCmhwqn0twv7LEyyJWfjMEC9D4I1x7gIuF/bbe
B6iwSRXSn6EkBbzI9j3M3cipKK1twsXiPlrJGBshGx8/9dn9qper5MfEC7EaNydZ
eBbqZAX+gYcMb92yhQVTppZi7bKnDmJk2L7CU1caK7KP8Swg9vjFGcS8YlbWbyai
SYkai46dOy0JV3pHKzbBlu7bCtUStPPY084GVOY/id1hY7O8+kGUGjkekRVBgY8s
F+jTnkEqsYOWZAaMlF6GcyQlQ71VIDqEQ0X1M52nsEq3RxAURDmRrzqKjVufprGs
jRyimDNAA7IKKrDJ2LPx+ehZNIZiMODqA0ziSrgEHZesSr7Zui9t8lpwz0/nMbXF
bpcD1FHXQt7thAiVdmFqY79rgRCBJBclmOzbXJvjz5QAtb9ghQnJZSJlkYJTUmsb
+kcxAHohzupu3a6QKYr3HMECy5qtErFr5PKeb/oFP/nIgowA76bzYybM3Lqh2V4N
prRkGMc0JZ4wmHExy8DZbAxj7b0ObiRh0z7yb/Zi5EeyWb/OH4OK2I5SzxsJC7/6
niXxCRZzypBRsbOd7mvPTbSUMezLgot28sfppFqB8cEUb9VMvc++ar8Y/2teIiHO
L95KL4EB/Jjo3zMDnV8f0IE8rV3tyx8xbhBmXsY0tauPtkX0Eox4SUtt3vbN9uPN
mAGjdHs48cq0pjdQugMArIX/N/eW1XVec7X6MAIAwBl4sOFJNOlNJDsfBXxh4itO
n/z5ATtKXGhYK3NV3ioW/B5NwOjaE/RX/y9CNi6k7ZJgKzYh9m7UOwU0bSZnuUY2
a5mEGosYPK6JbQoQs1smLl7DbgrKi2iNavdu+1OQcHB1fDBPNSmdSX8/nFKq8XC2
27nPB/m1gDq47HmtxFebiX2z1/IEjjvG6wXlTi9z352tlmWVgYXPtSNlf3zKtkwl
x+EyHuva63ayCSYd2hIYWI0pE/8xYFKibkiMvBqgDe++ur5qH5elURmR9/gE4ZER
QHcACipjrCnQccBagLfgT+oqi/QVDntZQS+6nZ1hIS9iQ4Fwfb/UM3JeHWbwZ3wu
6rUShWUFs723cxJ5oEX+QWjHrrbBWDM/R2Thyv0RBa7PDwdX1FnmEvIwbfjIbU5/
6nIiQpiiQ96xE3QxiWZTOtvn0lfUyZ1i61FdPA/wWb8D+Eu0PZXAv1MYNXGaBTKc
o66r7owpyvbXMYZqIRwD/cz4Du9i41LH4ijuC9LL3H7JsUafgxAoDOwdFCLcsIPv
oILi3wESmGJtCzCqS9vPocvDLU3I0Uxe0Rv71QqOKSvaJ3QxFxxwAPC/CNl3lo/i
/NZpltUBJzZ1nXIjfZlSclNichapUkADbmmS8pW2gAVuiMqnjrevOjxS6FpkokxT
OqFXTpLJ+z4rgJQSS79BssqPnQD86DeY18mKh7hEOZr4s30F6wc9vSCFA2y0Y+vF
wGbF8z5vaQ6D5sLrFKeFqJxv1sYyGs3xbuo3JgYX4qmtZi5eLi+XVPiTorpQdASE
vj2cLR93338IKF7KgAy0V8ariAoxo9bg6ObuwwXcSbjjRTriszbBxW4Mq7tNntHf
/TfeJIiHbI2pEfxO6WT3wNy1AI9LwlixJLDE2WZ2QV/Kz/g14SHA39fpAqgdmb+J
H33B3tBloCx9eCCuqnHqQhmu4m41NHTf7jjN/EN1zn06rsT7ZAvBqB486d2Pqre9
jUekpg91yfmnDh7bcMUpDAqEAc1Y1D8jrH13nNgdxnqPp8q0zUR+mMhyWLiCMEP0
RbmOTMgP/yEsFobK5D4dSrmknyhHrLwkr1klh5gWMK+Lx6vb2JN9NypKokYbPqrr
opLSoTKtHL6xRcpNV6uVXmtxMuzV5PdY2WLSobO4EOLJzzz+nG6E2B6+Zkolrh0B
08aGtIpDOyYLXefMKLK9tFtkh69hAo8bxEfkMYl+lcCBwMUAfj/TlueLwXgoSOh6
ZngsT/T3rXpxwqf6tukQ2Gsk3uyCwTZHn7lG0FArZjpJi+ztYMkRxBkGmvjJeaYW
JQUoqwzYpqQ7P5UoRFn4e9oezKZFiw1wVDJ4kkp4osit7GzXPJ6m9/c8Cezw8Wrt
d5Nld2btaKlYVhJ/4JYKu/bWjZjd+cOtqXJtLUJK2y7I9KjrZjqhFlvRnMWiG/Gr
63LMX1ZzxMp4V9NFw5tM1Zculxohmuq8tc9wkc8zM4s7/hiSUOClnHHvRZSHQ9Cu
CjXUEv31rlcuSCAxCkaQkp+yvkMsLCywVhWsZo+RZWELvL8DxhJU5GHCxI36+s3g
ks5yVv/HROmTMSElAcec18Vp40sLcORCd1DGBfGRjzsgQFITSaoyAo30COkeiX5P
VbVimeUdIXCWi9O03yOKo1PBWCufj5T7IlHpF0a/LX9aqw/TAFN8Ol8dL+9w7MmQ
/KpyZ/+9Vhh1KPd8Jk19eTULXoX4yB43LPXZskfjfvaXoVc1RBlzFB8iWuDXgC5p
2E0o+STMc/K7LVnNF7X0XNIc06ehZy5eRwxwNOsNoqzNS8FvXR/vdjwjUAkvT75O
IvBGCX2oWci85mFkk4Lhoe9p8cE5LOF52unu9TRSqximREu2b2QG/UPXAlpCxmml
sjCUwg0icJWPzsMYJU4ete+Q7rNWKJ6eeZIQHpcC2SpK6OGMgQ4xZDprbMO53eJ0
zM+/MGJDTLkHaOkBRpnhKh+aifIZHWrkmsxjyAFZQZ2YZ1LN+13CgpP5zFqkJRyC
C4+Qgi9Q+rDMRT+oEAdcUjlEBzi0TFij0HR+x+bbtvVngXRZvQCRntlQVQwiZwr6
UzCC+3Z+mFBYRkIs6YTcPj/JRe12e6AYgEFFxCbI4D99Q3fy5FqJQU++LAGANouw
Bvnvna6AefgaKRRCgU1Ja/xQ0MqhM3iN9ChNZv47v7yQV093sdm5L66vlpXiRudu
jf9+H+6D4jMq4AqAULi1oh2C6QJnrzlvQT41n7ZIgsTQRmAVB89lQgHQ/cUjQtBE
NxtgVDLHLppfOGCH9Y7ttNmt8hFiLs51LCFWZQYzF4xb6KlKoZDZS4iAAHK4xw5H
bN5aCW6E42IyXNIxdgkowzDfclQ7Hj5QwXRaodM3rtUOiiO1Zr8MNbPhMZp5yU3f
vqWpE8ysBsdZnh8jeqmBxDQuuxOsHfJiv7ggX4KNBpWPUSAqLbz5OnrNfPq1FMSC
jvbZKotrzbCd9ATXvcQHa57sY0fm7OZ3vBRnU79GkfYRnMNCFeEta/RfZFsd2md0
4WPQEj1Q1AaAsKqW+fs4py2HjySB/pyKgqCRYxrL1x7WITex5O1CldExYZfVHLn/
d2rioxlhPJ0uzMFjAWuX4DsRk9wFN1L3bGLJ31v+cfPNlvUX/g6or0HuRNjpZ/SJ
xICBaEMVWvZ6xfgUc8Z1uw6XtMs1RU4J6H9s4dhEPcBD6Xl4N2THFfO8wQMO2eix
aGyfAjMbEYabpH36vxvNLEssENAEvMPWoZuW4ov7hgX3BOlQeSm6tcK8Xfam5e7+
B/g0bBqUJrr1Kl2HA0sx/QTfFqkY0e+Hbj0FHNDHAUDRkiSt4iVHbXN1LvVwNq4N
3l3ZAouk0se0VP4GTFC+oyf/yL5kzAlVo9C8K+9iWbsqaQm1XIm4v39QC01i9u5N
MAhOwm9OcN+659FIF8W9zNS6LfH0D0HM38t1qLevp7ATGmGMylZUJKwP8MLpbHoH
goDCv8i8XfVSRqm521rPodZ02WxXJucm4o1untumwue53/qYdNatEeLcSYZly5Bf
H5n4rjwsR3xeWowe8Dg++QOztY+F5bUJjaMt4vZoU+j/ppzBKR+WC41L/VolUBC7
IvREDV1aXds7S1kmLffLPCG7Psns8IC/9o5Bib3M+ABj14V2Izy/YzLK9CjS6Qj4
YyAurGt2WlAWRrcBIF4K8TDbTSXp8iUYR3Wsk4jB+QMvoU+xv9Siq/BK0q88SErr
+opxeXqJ3HTvtUqXzJV1HcAKkjroJVE0F/s3sHM0G/OT2zsIhLHrj+Op+7STtg6S
3U5/uRm8vIvZt81Fn4QzQFXpHZm2uPVjLsVp1444Butgq+HWJTRnjNRblPpDcpiz
A69LZ8MBQKFjYosPhImfcrZr9LF/yTxGsO7XF5MKiWSSMRiSfOsgEg5vi113k63X
nMlzx1Io6g/bIktF82Ap+IWyVVkTuGLVfoJVcOtqvh7Fs+r6FioL6Fb3sN05pLer
WMHsOnGEzyqwJtFqw53J4v5rxOAOM6xCfEuMWiJT7Yng87Rp2r6HPgElfAqRo6hO
lRZE1JQ6oM0VThr3XH3eaUarpgT09t9LjI8BNjVfQ+hMPGo65t+cMyjvpWYboWkR
Nj7akg5Xbi9Nij6MOUpbIbnQZu9e7mCZA8qV1OGJljc8KDStmslIA1vB7zzpBX8d
6/Wc8htiBrQ1qap056jYx0ea1ChqP2lNniXh+Q6YORkQYVsW4nuFpI68JtrtlsnS
8SaDfrvMkJ5Z4IPluloX3GkAyhiKpIRsNi8zn3YweOjoE7ctEEqgLTq81XkVb7t2
ahyhCzs1hjRLwt6qwfL7Qo3MakplH8GwI+5BxyysR9mmuKMgZUPyH0uVt7OBBNvD
61Ub/249lyxghcu50q5TFufIqxDaUjniMj2XsphgPeD68n9vv0QO7LDpjm+dRMth
M574NbIh3lCjbamq2XuSkNmloplLtYrLPMIMsxGOx4c7CXLmAV5RYwMDuelv78Aj
baQF21v4JyFFw4JU9exwcW+DfpzPE6KuNqO/XJnTj9pov/2xgYqgDmKlEKNBTFlx
mXGDieF7S9Ggxb/2+YX2Cf3Z/iO2qMg7fGYTqoRVo0VaRsnjKux1l7zjb6U0TceT
9XEu+t9T8vxxD6nuFwefbNn3JWkiCtFLJrXQXcDDEIFcITSoPzvV64cV3/xRi7Sy
X40MW0qhBSCqR7suW5UJTGIi5b7Ggzpw4tuq6MRFQiDE5e0WLrcyxWRmrL289xn3
dLKJ3PxBeCPCnfwXpaF1jiPPTVyqRlRr1DPw9OarFo1JfXQpPvtDp/pg0EoEtoHF
FJlRhgoD1XGbQHc56yg/psrNYDZzXWUvr4r3Rsx+/eCDC9U8PIqwAJ/IjvcLLGtZ
5se3TojAb8EoqP+54WpA07J/hc+r6AEX1f6Oluci5O0RlFqBwXneQIs5hAx68Ggf
YmJzMAWH9gNJUrx7Y3wEIpU1kDRMGXeV///9rLA/keymS8GntP1ASmEESas2PaAK
Ak8k6bNvy3YK/opd/uiBAJSHqjFwYvrICrjYHoppFfVx2r/ceUzsuHC5pi+MTRUO
+cWK3CkURQQMkwskALltaWDx3XyZT4FMqbHvjSHEsDzXmlknIM8QmanaEiIfmcI1
fegIQPOkap7l8IRdGX8hDFdL2R7jT+Bu7AYYZydzCgx+AIy/oFoYWh0Q1X8laTe2
FuURlyXx+w5HmCKODoDDTsC91z2M/BfYWBuXpuXkJ/xp/DAo1torDDljhPg8CsE8
2IbZ7PYh2GD+E8Pt5mR1Xvf/s2Aah5mKeMPSHbE2LBnDCDYKW2F3RQMlD80yL0fV
HVhf5kfBmCz8MfRLZRoD3WQnwzaDcIsHWRcu0MbSnktSBA9PZA4jgJKp1+iJiBm/
VmS9Qf1nGYnvKv+VwOgjRFzLe4GmAYGS9N8DAUHJQvepErvDYd4gZCoCUk2ElSA4
DgGFANMsaiiKlpEqRY5yTH79MWPoUjSu3CxuSUWwadUXYgn9UyCFOGH46o4Sz+wQ
kZ+aE6vCJGlM6hAWMvcKX3C2/HDE9Zz0hfTFwEf/WYFn+etNXa0TRe8Wb1PKRG3/
g2rmvHOQ0VvRvEyn2+CkzWiuB/UNr5l0xXZkHKcruaoveuOHdvOw+mVyiX1Ic8vb
n2xChXFLhuFGcEkffD9mZ/NOvxXQ8qXqkTuZOt11UhiUfVLMwnAjjZ8+Y4Ctk0Kk
LOg7iK16GjNSTrr3ngVo3pYY0He+uF5aY7M1neVLdH1vWfmTsbjUEhzaIlCyBlnd
SaA3heG+IFfqzTAGvL9zzDQH7S4bkztwLzX+8LP+cr4XkIi7vYG24nsf0xlxmspl
rJv2YtKgyyvPWT+CIcEsgDG/NocA27p5Fani/VVyg7hXETffjDikJpjnqBGHCHVj
vigq3f6tEzSiOR2SZxr2kjlcog5GWeptRhrFfkPRXeGpjUQSNnpCQebBsxVKz+5j
K44+4Yf6dkNGWLR77hOXKw6eORDTASuYMnbDEdK2jZ7Z1d7Elguk8W/QUovCizUv
/gitF9Sx2hXTTuIjjhLwhstN6uaD4QVl7SWlnANmwS3j1jNuVbH3MLe+OawQW8Ok
7SfuQaJCG8POp1nkLsBm563Vssgq2oB8u9QhJ/fMatRQ/gDkQCuXAKNZYKhltPmt
bGT8Ir/mV3TfFfy1+ZXDHnnhZ6OyUXkLNELC89iDlFK5ivsCiNqUaAHmD4yfb6fV
ujur5w6S20Xdi0WoKS8+mYgollbjIsAvsklfQEUWiyuJ5ht9y1yx3kO1TN5Dd5iA
qHSMkjXCQEys/sHHs60SlSmTQ9MjpCjxrJpK38lCNFkzODYOJbCh46NvzhKaTvyS
mVCutEZg2Rbg5Fak9h9PtYfuDPsppxyZ5BRZebUjDh1CL/iIAz+v5khuWffkxflD
r+ts8ltYlqWceOr3g4FCGcCFT8Fdd4XoIKTVbPhSoB/LCMfjGlCQhvzDVM5zdsU4
/6TbIXdtWqu9wiPfPhU60ldmvtI/wkeQ1DCpVp6gt3or/JoNZvHmdfw5KUlCN/2G
AGqOBdiGG7uUlAwifqHB7pyKGmMRISkhrEFU8XyptdWCsEN+QL2jLysXcJ8XsqYe
1PNrxGe6QwFnFEHue431ExNzDDM0So4k2kPQ0v2eR5lUnhhs1U9R3dmdIuXt21E2
ZqxYSsUD1I8KjZjOEWTcYs8wD4DM8KOdC7j4e4E/PRASEc87iA1bx9ORdsu//p3P
RsdXG66tFaMjTOAvuiCzx83XO0rugWxn5kXNn4M0x6Btzmjw5zAg9/oYaQALAVg/
z7614tXDRbEh34+7C/6xzCAThr1iWyyZ1spC9PWrIXGK4tIcBkCK/fWopqUfxktD
UckFN1kjV/3KGr+sGF3hjWNnkKuum1Uh1b3FqLCmmDfIhCstlRN6WdkkrrUL5aj9
iL3d7y6tGv4Qce44kPECLxlctDF8bJcoNBBJXIapQPpjBh+V0UsnWNOMjBsbLg6j
n4XWw9foZm9yjFJzsxdeLk5qlMQ5K8wO5CE3sNlS5tvlHa0Zm0/mGi3KGkKdInsz
TRovMtJ9RsODEPEYtK/fGaNrM9zrY4UQRrxNSHssKZXCiE7x60s4hQZKv6bvFI2p
t/MJjkGbATh9JIIMzki6KKoi/N9e7qVLTqKeOCr6i6c7FJGOPgh+y4oYszFdAzN7
HBGX2WMiixmTwrx4mR3GFdkGN9X4xaTalvdfdN0aVOLk1ozsdo7WyvAmnaALgB4P
gUnEuUut8+ZhZVwkEkag74eChPdRVDubRVo4mSeb9OeLKIRKKPUOjO4zvLmuE5QQ
pRQV+nEXeFw3VJy+HZvLdadTlhxJuOzQ5cD6DJoOwpHtbI2x6FxXtWS8eI2Zjq1y
i1+pGeyVbcEx4MmeQINQPRXELFfNGm+GqrlmHKS2Hzy/qLQtpgFAegpEBoqgcn0z
4UcDjGv7Srbl5KtAnbdMfn4bJ/DWmoaXNhpA/89tavVn3YBVB2DmG4v9qy088Mjy
qPP/tMJ1UC239zGZXpQiJrCSDLPyuKcewIbuz8e7N4Yviw1sqJ7s7qACrDodEB4i
UL20/flj1IXh2PYs822kC8zx89y80tMFLTjGsv/106qmOjdAjGrVN6Uz+KxSTn/3
e4DzAKSNZxM+oofCvHKu3ittJGjlip9SAE9EvwJuns9q2hgzJjuaYfbiU3TDoLI9
1jCIdFEAfRGe3ZmUqZtFJpmwyPKxANWOUeN8wZsah0QXGsSaJLii40Hkti1cZIC4
lycdC8d800V8gy9L1IBJasuCHVSfkVKNlpBSR18SXEvA1JY/rZeOh28mrxyrTqyh
riuxYBElLanAqVHXsrmo6X1KaeafdtE0M3BHDfpIzK7yNghN2hTkyHmBxzPFAzqJ
ofR5FLvE9GZYxA3t0w+1zV+r1HD/CoWMZg9LsNRAkBCaU7/BT6uE3+wJ7NtpXIUF
eptIPg+caRiwPUX2LIxZggJqF2rmP2knHWFixncEZ4coPGBUtHDECtXZrdrMR6Yv
+42rMR1Xg3GCwlMC5KgiLixpmQTCOjOzEI3cOGNBNX0KYaRAOZxGEF3q+LrLsGW6
b5F2O9mTi3UWiv0cTc42POEHlEM+FudUpmDxU8PkxvTsL2KYDqu1x6dMI6+6z7Rh
A51vRdNXbSjz4Iieyq9oCMOqqrmXk7q8f59KXBPUY1DdTWRnq+h1yXies3NV+/ON
AHJDwwCukIBMPGirNIr9HHDLMLAMW0fXDZkce7mv9bMtGKbCQzZNrQ/JQiWLDnfG
H/SJOXTTyUrCj9LKhuFLXQ7qxofQKAY+YlTRepBYqz8fBzPsSEdW1lxmXTGiVhF8
NE4KWqpOxMXKdK5HjX/er/mLOAyiwUOTr9tPtTI2OFrZ31CB23KvpahyDl6GYA9E
oSpgupSyQWkeii86vmhBdwxlOQlmCJ73a9vguhPb2cxXNXz6caLHCrGduQS8jeHR
JbtlE1VjBW1LrFQr616jrbkcoyCXJyOyAq0UGMMs7ITmlD89bDiwtBegM6bV1lzU
glL/OWSrGueegZz34Oc5jRrs51Da+ytK5H4EQxAj38OPu/gdJXVkSjJJ5mJBDOw2
X0lf4G07xrenzKAFfWv7C10dKvC21hATwNkpRqo0eNB//9DKlh9JjBIJpfe8wrBm
dJxr9TQwM0nhYAQxx6x87583gXnQJgOWiLirwjA04gP1nFMW82xP+dOstwEMappm
dqneKJtmT3IJm0Hasvwso15TZvcSoG4lnbnVIUqxCiWiyH/5SsFpdAfLdb3K9xUj
BcueMbGM2ChZsDFyb647NuhKJzsqArLNX029kd1pdZspHM1CShXUahOvf9LH70PW
EJYHvpGyLLOeivhO/K7wAgIaO1VFXNRD/Xj5AAqXZjVJQtwpmvvmFDWMztAWynj7
6bJv+/gXYN8lvB1sQoqVuk8yRSBVlFe6IjvLtS9+YJpinL9DWVhAOoy4c1oJWzEe
pT56i6rfFy01KKmKN+hp4fJ/Q8dKYOGs8DgOWBdM7mA9lzc5VMWlgy7cqf5SoKEf
Phjz1Tk2mAaeIncMxdy1IHwMedpEYTjLmiDaOrqrMUwkDf3wNznIz5bd9yd7V6FV
WArq1GspAVdBllR4OUzB2ZVR+RUCgAKmusqNhUIba9RxIXfe0RjGS5ubasQDFKcA
qfcr5Z4qYtMA67dYEhR6GhV0TyBylexQovF/Cy9ZdxRh00ju4mUyOq7Zfw+Vhd/w
BAHxsxv7kGQ2+kxKMIUzvb/6CUnxHZUbgCEKHfWyT3DObasSuc0NY0F/4BT8uVGy
Dy/vQoiE+POLx4Ds5Lb7EWTmCKJRU7/wyWuK81HCj+WOPt3LAf3d7LnZP4A6sXRk
w7MAkmabiJFqcRNP6eCrQNrlxCIg5TgphCQx4MoNzyL6Hu5M9NpVwLbuK2M1iHV6
U2YboXFdikyv+Qtgp+33OKhLUkkmrmjv+NA7zRL97ln8QSgBBs/2RGkghi8aC4Vc
hYcvSbbmw62jvbw4d6iY6FY8TiBQi68ay/inS+cDMxI0U7JRfPQ4ZevFCShb4Ikl
p8fhx1OBBhKAhp3ukqfxeBhZtpjWJrbZ9E6sk5DNlMEIGaUqvq8E1Dqhvb8bGSGz
UfT5SNUo50+Qc59/rPIAyUpFF3k1mb/lA79OyVw4rANeJlSsncry2iv4QxTGNAiH
QBWmbaLOahJl6e3//p8esPEBFYFF19E+Rda+7DSrDv5ExQvDuAvz9Y7+4sr9xQHD
TxGmiCDFCkhn06I1zd3zpFk/lze2oaHrnVOZFfpNgge/T3FtFOLJ4UWltlWlZVsS
9/6NoLyb/QdfacloQJduuq3lP8IKyHSFRBQ6vBlqnFy/KAqWMBDaFJ1BsalpuT8M
Pk1SxV7B7g44INyKCThNpsfFXvn6mTI4GmRkFrQpP10lUr/a9lm/K/DM7wzdIsmu
yMHi9IQctPXSaQZ4pMOBDOItdEXb3Svi1M3QbDCh9yR5bbZIRUTmGvPukiOqHXhk
SxzXy5Ca7jyw3HmMRM0COuMphjzfX6PhGMXVEYIBU+jmZVoHp87CoduGQH4XSvjU
mzxoE/WiX0+akwIUDp/1scSZET5TR+8YXzhzz3JJpB5t98LTolGgb9Vlu+rYjPPl
UJ30kIdxkIt1Ybt5dzK4ANTeA3SKkXeZ9n0mj94DX6nqoLalZ7eqjesis6/z6RJc
kFneiAnvtHF80+WzHsNozGdiQfteo9dQMa5KYG98sCVG2uN7xAiyPJlXFd8vrviD
sRbRR03xWBLjlAzGhsByDC7whj2SdcOIuobLf7RnplpgcfFjnrJjO041iegeOItF
sFKFy6Yxwex0Wc1EghnMlTiAMXKmrt8bJKZCyqEUDLX4tgtCDqHPMcb6yRlKeTcf
eAYV0IlvNXa6D5wTPpgtfbreN7L21LJoKdhDbmXmQ+dHTGJreDHkBwOjPAh8xNc1
05+8TIXvOUN0y/X5nTLsYNkBdycUAhV6u/h8NgVQRPDSm6il1bDBWQaQwhRnPkdY
rZdz521QLOlLQKqgh5WjERE5ssmhPk+7alcdPaI+nq3MaZMN324QvOUzcBnJQzAm
cdljpATgohit+SOVVRzB6S+xySupMvg5FqwbamMlt2FnZDxLkQbPDx2cO6weh+Q7
VhMhrCeszrHycDUjjPgp2I7EzrdVg+yqDOrikBgQCV87vKmlRDIDBsOcBIA2gJJg
E5gkwIncet2xtrFRgrgxCmvR9RpkVyJdCFpQVIScMmyNTOPrtgiQTXSu86YBZv3U
fk8jqyNjQPa1fwc7foE1nXeZa1clhGoHbIzme5/N13h7adaiDtMMJFC0VmI7jj9Y
0s1vC6Ha5EJgYuWTX0v4LQHw8603V35k3p7YwXSZk0MRPfoXZeZ3PvZQ+mB+6yhQ
E6W8NPAmBtuMsXPjujS/d+T527nQT5vF0G54VuSqADJfvG5/HubiKiZ8He/gx/+q
CMcwygszrTGzreyg3LMpEq2QVpUUK/PtqB8pgmiLbzqw4YHBsp1jOGO9IfNtXV4E
C7Yq4M84dsjYczVcdQ2PdFNji51v+eF1oV5aWOjR/Uon6DvZwrY/tK+c8yUQdN9O
iRyw/ckX0+B3WtrvY/rxpxjLSnwy/47RgbOGIJ73INVbeEi44oigv4oPsapwGXNs
dOqpMlJuVLHMQabCna6lBvOw2vDrqpjondeGu1WcARPSup0TPFjoGzAsoS6Vv6g1
9RZoD7wPpM4C2Hg7f8aDANzL0B07YfvtWwYXG/NaSQy8NYLR0fm4oFHMI43e/6rL
nMHtVev/CzweryajH0Yv6AKqVH16cv1A7FR30NjkoKGCkSLymGr1u+fUuxc5NSJG
EhW9dUC7Icb+sXXBZA7pwSwfAlXesYc+//paE0tMAxzh/YdSEnQRPnHe4pKVonkP
x+AIr8LLrs8rb575h0c9kihmTR8dI7ODVNH2rZXGo/ul73H3QaLgpTxtxAu76ZR+
ag9RcdZnyjW34OxrHsvPlPpXonBsLWwlw49XVQrkuB8DforiWfDHj2FydWAEKTby
+irH6CENOjghHmc/0bc7HzYnoeUJYrfGMvb7oTi1mY8vldSpOOnD5zB6KrF18YLe
yz4V189mk+caCLxr+/RRd7/Ikz8uRcPCSBmP6Uub9f5PyI5xongdMJRKGs4d3uor
KslRAg68WXtUbxtjhP4YUrQE5skj7db/a5r1huSiD3HSLoNQe7HxhSDhplg95tNf
B5kiGdhzvsZx+QedQXY1Vd2uRB3sJ7W8RLzj3Cqn2ePgvx/8Gv6wiR7HcGg8VMYd
7UYwGtoYMy7NyU3nwrPYb8+vCXrhkKPfInWNen8M639UX0pPCj3bak3KZNJENbjW
VUWwXY3ZYZOo9EgXong+7eO4jThhHsRwtENGobP+04jnM9s6LK8GuRVstmTh/AmV
21PtRflWzAsd+jT6giCx+9S8iyWhWnYRODqV2GUueu0rUTz9WHOW24v02lRl6uYg
H/PfUspjYk5pjzLCpmpqtucsF8vkfsBC7/3lFgr5uwu4Kdfg6g/WKkG4EGaJEmDV
N/I01rWRO8N123QnFJny6YjgUOsnPdTF/3sZS1ekStmaVjc/gSYC0ToKK2ZfULaC
xdOV9De8NCZHBgjBq+2+fk0VpPpDH7imjYNMctq1oEbdNjkWp/E1cecjxPKpL3ZA
PryMdJmzNhnLsuCYTExJpfFG8gIWlQ0JW4HP4pm7uRFZhJd8msxSgfCFc5TIn0iN
OaU3BMVhRppI2gvAZ64rZK8uK5AnpinOY5Te82Oof8mGQpeh6zc4HTFf7AkNkVYf
Ivn8C0VOevgYMs78Mzvz0qfpbuuehtb/PC51KJJYBWOwNfyHRy1Ri9Ocbarttlz8
e4+eLdht3xaD5VsL8rx61d8LBfbXgJrmedFJgmJKDk9hNeTTNZxwRcwSSb6eRpiW
fejLwaHILNjMiZeAEQG4vceb5Y4V56pJER4OXS/ssjwdhFNn5A6bdeFZ9L+Khua5
N2uG1bF4Gke14KJWxtIKY4gfnRzlZaCv3w/zUBQAhS7ENG2AUljsdmlmkn4SrKJz
uS2LBQCzPeLJ81z7Mp+tVWLfFu9SXZWSnvBTuOHDe3vJFK/vgMEcfYR6mNyZtAWd
zGnnUXIBWkU01ynbz7G7PVkyP7sibBesOp/zau32vTYRtWQ+sKsAXgrsTKmz4Vs/
Uv5aL5NfJRsL1/RweKwgoiDF2TA66ByI3OeJcO1PfPk0CGanIMjDIcnqaSm7Rgyc
AO9kM1eIvaJ006+ayuv283i6uzcKgJ19pVWwIbs2RovgjwqYWAA1pFv+HWbokW7b
cDxFA7NXVL3wO90ARIBzI+82GsJ9qT0xqWriJcNX+Fl/IIaKn9rfTfrim3HtwLbG
PSWY/uWCK+3/506Ci+3pwdXru+Mp9mBrLrSjpR7MbMvXEQAbLMi7rkZC1sKK/ZSu
d6zvE2QiKmdF8Z5uyDNikzOcBwdMZMAWFScuze9YvecNACL/VbmgzFbAaFYOaW77
D+1gvJ7bJXvZQaOlDIT8MBbUfWae1tFuIojIU5sHvmo+9J1jQgt5fO5VEpGxjivI
BWEKjg8k1HefvTexyCZNmc7qY9vtHMUjvvqCQ1BgqUtIatKhsaxK+Ythw3QTlWhd
cwpoZXkaDAAFe6V8b5BZNt6sjZuV67UNJYt55mGo874hMNCutW1AR4ZVQk9DJ+Cg
LVx5nGGKh9lWFk2HiXFGzUvYSLi/hNxG+0h+8ResueYGPTVr1jeypj37IGvLezO+
LeBsfY9U+gXZmvHvkrvg7QLz/GjtIkQ24XPvNGxYe0/LSdSgjqBPxPSBucP9QVcg
0ZqzOygRcEuVKwXoFStmruUZjRwDWWSv8j+GkUxOz9IpOQB3S0qiwpKZnnO7Ntvc
peYbLgrR5qGnvgATKJqR2pd8zfaDWlNK2GM53jU0TVNlw7/etibSffFglZkfupEE
TzisargYQr8mO5UgnxHwromf2x/g7S4Gqd9Hy8MFac95uImWTYHzrFQoiCE648Wh
0iMq9YydhipiIBLvn8lTMjposJofscn7COnq6ZRSUUY7a3tYh0Pn+kVBA/etqFUT
Ebe951gxWaddRc1IoeIAnO51l7Pw5ymauhbp1L11kccPu8+0NCFwSeHOMESdwFu9
iWxixfuOQAkRAQDwcF+QR4NmKxMkfkaunfCFJC8pppDSqj6H/ABrHR6OM5kiI7pQ
sjOSjeU/XsQuvOCXUE3Yb2+udhmGVp1bZ9YKwj5rAmInzTkCOHp3fQuOBi507vkT
K7AxoAr1/SKmfXLPACUGoRVVpvB736b/n8zqO1w4BAQC80gzuT5cRKM+kWS2gX1b
CamgL6BsAFzNg6LkyRbD0TDN1auiBqtK6n67SD+t9tQytvquPsdzTb+7SaTjnwfZ
JLktEDq4yQ6zfQ0DjGDa3o+J98RJStulEZBjxNQRxQbPDmwdnIWNmqRwzY074EHh
sKAuZUR+wV7x0rEbp50q8vpaGcCAeqyvozlOUxXbRfUv4yT7912MGyFjeUuDmo9O
rpD2IydwahDGYEPnoeS5Fo8L7xQmpd2v+6gNzslb4BJC+VL5WjCTwARS7lj6tW+e
I0+NqWpIQ6bLk2cASJPt4OqHHlonFf3kJgz0ft+Li0xquUuO69CQWf3AekkmRZ9X
cDwS2WrtFHhRv7OGPlXLqlKJGRl977SRRVJoXB4+DZUd/LZiyH4ovnMEDiSA4sLc
1pxUue3TYp4pMOlOE+EfA1ioyetX0d8kzJZXE1IbiW/gtYDNXCk5xwUjYejtNQf/
iXynXpVOFtT1NaR8xNg0XnJdhlSPA7wz4cj8I35c+l9X2PSA51KZXv5gnwRjNQPr
AJPieN1pSNJ8iwUphqdedqW/gUdl/i6Sy29NgF3jWnKwUdpNoOeCkurvdXf/8UuL
M2V0HboTW2B9yiwaPJogRjtyvSzFBGQrOrZLHs+uE0Br51KLY6JaX2Loa940NC9+
G/Uel9qjcQf8FCFSp6r5x2IjVO+3OvAmPfIbUsBWWQLRuWZbSYrKXghaTcUcDA7J
VLDYrLISbkUYCkR2ExD9ebREF9qKtKSNEikRrlrJwV6+LaIQczLpiz0g34xOVKk1
WEm4tUGJpqXfNbLNC9XlG2OBnwQWMDPrayhEZhXExWMD8VPAmEhZNcUtHmITtAYD
SXnBE6i4E+SK4FDjuuv3pcRwHFIi2XiVsEUE/nBUxFhLD3uHmKJSScYLzwdC4rAA
n2XHuXwCSC0c1T7ZQUW6dcN36V0yEf5IropaA32oN0WLRp8IfZ3VPX7KUn++a+NK
cbVj2LgaRZ7vZd3Fx6R9tyHgi7L7jkLEQFC2cS7h20pl2XsVpvlTojnO2vbbTFyC
1YVbypxPqAkx+7g/D3eH4C5tDrqilLxEMcEgidv7TFp86atL6Bq42NwiLIC3bC0v
D7Zh9D2s/thhro97RMdpgH7Ze2LYkTGqfpjUnPCd/hiMeJrSXrC/bCSwaDFXF4QD
AV9h4AZHQLJhBnmCoKhcdxxPBfhHe0yatjW7F8oS+AEWIXiKKL4rEUpdzCD75tEi
tq4scfkurOVdROZYjRlWQ0RG3t/HNF5kgUAlLMeGKS5kyiOp6jj8y69aI+Cwd4fM
A9e+eCCzCZUKoiYrspP9h5rF9/0jmeLG9923c1X4n3F7jAbMcRt0DPrOlmh5WyRs
Ks4IQS6aM/H/2EzaSeEvwgyXr1HpzR9T4oLVRRPt4HIC956K7PUmv3Mo/ljoWjuH
SIGewtSm7XDzX30Xp+1nZoJ0vYm5Df4juWCW79/jPvfeX3AfvKowbIUwp54YY2nk
QThQOKQCWnkZUZTpGFtnTTfT5bM+Ljt5Z5Rs2aa8lv+9STOXtcsVup76JZPwTB09
l5tmQruMPT242PLA9LlutC426BWR9j/NCZXfMRGQ0N6fWPhanR6OPnNXSkIdQK4b
dHhOfSGVK6SGECi+ceu0tvKaanOCFoTk2TbspCWmBD46Tv7vRb2yd8WhdcsYgWlI
AKswDylEi6pIa7v7yLfPpay4MNr0oFKcvQPmScb3YRoQfvxSXhHIWxF99ru16WL3
+H0v7sbOAE1ld/5Ypv/xu0qhHCk01dQ4TrsspotOuExqdvXl2UyxIsS9Bkk8KJn6
nSX/X+bhcySkUwIrUV3RzO7nSuA4TPOBr6RGt0XiGJEqw+3Zf0KlcYGQc/kwSKHV
8ZL5M/zgogATaAmr2WkuXUdRd1rRFSu31XrL7Ab5Ehw0mB/l+Ifw6vpnluvj4vVQ
2HWigmtVPl5PuLZlmieJzYFrLivABJe3EqmN+R9oOhi02mKIWQ2sw2P8D3M1u+bJ
ebVxqiqUe2DhLZ9EwLMnpWRYnOtVWwidCfrntP/AlbesArOHLtLnCWUk+S+vitCO
QMcua+oJ3eEBQAkQ+g7J8AY6FN6Cu+faboY2Fxp2kEBEvLa8UiuOmfnRkoP12k72
/U+jATEAy+nff59t8LDnP4IZWODJxJbPkf3hWwUoqmBNLTDA3tvOfLM1tWd3zqCO
GrN8S8aQyTp7fu2IY08MSn7c51a+3Y8hJ7sK8LIPU7Ln+LZChwYDvPtK0DNQqEkx
4RI1QPaSdydjhNGkdDIBisBkFNrWPffAFE8ITPtHQKOo+3MagY8tY07lqYtazyGi
SimuHJdJRjEA7XN7obNycLKCD3oBtuI4rS9RTvdgGuOXgrntAS1ga/TO73PEumeh
S6EUaGlGtn4C73RT9BcfiswX3AJskxCjEN51O2JubiB5comEdx0Y73tD3N/OSDmm
99jLnCmkZt0FrrBly10D3V+uBe0pJiLQ332Ih5HR6zgU86dtHoFSJaywD2KTwgYB
AZ+SimLHVwhGgXtTSP76gNpmIbkvRi5X3jIduw8NkZ/kA1aTE0IKCRMA97FmOi2g
ufy0NFGNRpa+BcUkstJfvxeJ30DDqG1bfDccozLLqj0qPM+k221wq9HzP0HAhqb8
s4AxvaSsGOnEWKDybPkKSZ464/PhaKYFepnskXbX7QfSOsKFUp3kfV5vah8Z+59J
88iNmh4TpZBEtoqotXks3f0WBumPYN7n8yIKoszdCFwrHMIaYWowvpQKCBDxVy1H
W/A2i+B2QUQNqJ0yLcF25mUZCyTi2aFzMij6KM3MzdhVSob0qo/qO2FTYGms/tm4
tj0j2JnT0pJzHTVGT0WTkTIVfCCosqn6fGLCdTzC+S5wfEQ82vFPOqeP28GjdCr8
NrWXbrc4t8hI6aL3olMZ/XkSoeeqs5sV5QjIcYZkBZezqHwH++Y1NAsXWp4ZjHNY
xFi6GZz0GvLUDdugoNBxNc9nSYYWOAuBwPaUwA7aq5c2OPDpCaZlpybtuZ0+p8jN
ljvoeEEppWv7qV6Kp0wYnhWCpZevdLkjluYCP0wAEJkzT22xkvzIwWy7o/GP7+gq
CI4qc8rI5gFnicYaFxIQ7uH74x3UhtFOuRi3QFo+9zjwbUsBCPkNY0BBrvbvaIfn
6yAI2u+0nqHb4FtPwuEOXpUYGobkBNIiq+Pz7hc45oW2FSOsONqd/nsDv30pp7uG
q7s2GRNZPFrfX4ALcQq6GlB186/9g8mwhYY5xeeL0ISOqTMmkpw/RAY95Z8LEphp
AOjvaBBV2svw93VPR55CbS70AwtE+xO1TY1Zy5S0QntIzbgbhYQIMu5b6PxolQNs
hwj2vzUffGJHtWHUiZZkUm1ftXwr9qd3VPZxCLfnRbqopDgmAnpCVFPyMenGfEB5
e3eTtTkcYYk2Sl8eSIDZVEB3K18+zy/Exo+AsVER5MYTX2RBhsXo0cR92bSwUgZ0
mee0iUCoLKMg3gAESe0Yjdg3ydmWx3aOaR8vrB5lE61v2L1dVMOmIGV21YBSFHF9
Y4sG33wGhOqIhdCUPEn/EcWoqDcJE8khH/Cefw/wGIfweYlDf+TzzPjJk/sMvT+n
DWrvmQ5uC7aDYxRmz3hjOu5PtrMvQ2NiqFPHSxtEBVO7QoqreDrdoBaL829eUnQ9
UfkqP1WofCC8/lnEiefiM4ghtDStvWmn66DBarLmLTvNs2qGhfLg5oUZoRlVrAfx
OtMteTQjLNnZ8SoHxO+fCi+jmdqFzl5wB5GaRi25eWHi+tCK5WWAtdkMqDB/4xZZ
p8aLHyShOTjEAfq9hI+p6n71Xs+/xJrEcYI5D3futJ1hc6s/pOIesrJ29Wp2sSZF
H2w8jlFiJWkr1RbSPvYniqPXoeynzt/Xl1atS4J7YPJzdF8ZNUSCacwe0d/jMT/I
NR7F0r0vuoJ4yWEnckk5K4xuWcVx1dHzEKKvEWbsvWzNRncibEv6vXrfzSZIBIgF
sPtOBRdVaeXB3Y9na2H6yix5xEvzafurz/68Dc3aj628z0NQdZZANG9kp/GWMYRW
zS2XDv5w9qujo52bXV5ILA5HPX6G9JkDKj2Liu3Jlams7bwUEkC6/uuAV6PMFv2Z
Fbrx8lsKXOmcd70M7O7NE3KWMBblhTHS3zj89PRy8Y9Fa2EwV0cXN0qk69EOeCzo
Pcu1SeNaqXQRzR19hPp1ixyRz+wQgSogZiTGN7W/JrZ0aRR6s+gSJVgF7hFxmNk/
cw/57Fn9/fcl0RwJigLJ+9HLXuCOA2PszlE55adsq+K7XlIgiOw/2JON/4FjTC1f
VHiccpBbb3SSrdgNPE2dZsRH+IxPAPHNftH/s27XK5V9P3KmIjBghk0SMXJnsqOF
KWRn/zSAmRDrLqJvabKpAaKtLINsYz89EiOCpSHCZ8ViJA2EM2a5N8Mib+rrDuXM
+1JuNo4lqRhEis9ymJoulR2L6S+Hz4sloeDJmyhS6ViL5foSp5+5AaRAllAEpkcj
/Z6JRgzUCiTt4JbpO10OFZPsvstcbRswoVS+TJn3brLqG84HYUyg7iZX1TfjwcNj
YuJZtoiyXKaPxTxUwRl4PrzngME6lRYmEhUdJDwML1knc+TYPJb3/4XPGYPqSaKw
jrvjeGQ/rNIa77nb8gLPD6zpKTkkG2p1EUKDPSu5rSp/EfJbrHByXKvSMaRBY6iz
6K2MSbxADW1GpzDy2iaMKkKi/aY34XhVDp+y418sqnNZqnKjxVJR/nDKRVZHd5Fx
Dw6sisKd67QPavgPSAi8tH85DUQ5La/Vemx18Pz+ga1McOApBermnZJwD9b5NBif
AqE/GzO7OY3rcQ6JtZcjiyCZWTX+5GqhZJaKw/GGZjD7PmROwePOhxN3rtn6ddOe
1Gp2MCqwis0go9ymCAMg8+d7E41mUvdVe2vvwWujoSVDQdmn8vzgoUs9UL+/Cykj
IPVSR+ykZxXERFSZdx/9d3aS9z6IObwyXBoiHuSalm/uAUqJE2B2i+iD81MONSgq
chJbmMOALOsT66jXk047BIW3BAX5Vk2A+KJKChAAbESfbGMqaw2vnslID58YXGgG
rl5O/troLYhNzqzBWYRXr86gCXv0Meyyp7q0bex59y0OdJekKQriIerlRj9S2PUq
aladdMGzjFf6AtERLdI0iknRZE5qOJqaT2IUHX8bLBvTzpjRWv+wNRyPneF6/DL0
xegCzi9/eQ4Nuby2Xl8M1obtMVEzglJg+3PGwWjkFdCAEuoTGj/BoedDpqGxI2DF
IjGRzLxOFM99sh6m1UOYhezQxcwkTZPw1HTjydD52O/9k8KrqKCKAaJ/7lTdCMfe
0vhfqE8d1/m+35QFAn7zDqzRTOZlKd6hGVgM5t8MNqd0MywvbFwbcWcvdjR+/3dW
lkzyjDQSGzYPyo/8gVNS1yfjrP6L8TUc59fsloypegWC/4X45BBzfrT9+UA2oVeG
KPjnyOdeVSmwZU/+UZHfmc/f3LK9UX0EJbeZbTPXW4AcPfNz67/yd4qC/qMoXnJ+
g89CcNqQ+a08m41kFhHc4LZS5DdMQJlGPgRNXGjiUCAu+PEOjOsDiJB9AWGTfNWZ
OCS3kQoPxU4n2qss+VQXvI5SwRFd+Qk/yt1VLfx8tZW+RbCev3NvIx+SyMCclWcg
ZYbmwjcbr3k4B19UKUJlUtfVNc/unUMpfrPHov2oQ6KHA7AiiOHw7w2wIn5uj5db
kJuMkmR8ZLL5qPIuCeYJwzbBiNofG5b/EyN6SQPB3dJBIc13fHRcpfE0hEzpK6gq
RWERFCqmodH9pl5tuiImFgQFiXIbMBmdLKMlnM6BPBBp9d6BcHzX9X9dxaZx8nCk
xZV/WfNLIKDcQUO2q9tpntBeUVav2Tj5bLgjtZQhRGfbm8+664w9vDjOIlC1xNjG
X6uxqv5Dut7W3AfzU4S8G2BCBJ2muXNa/ngnl24i/exJfqq0K6V6/yYEo4VR0Zlq
mpSH83SDuZWvV66D61DEMFTf4N1YhKdiOVTSiTUPFNeEyhf36nTxomFNwQuvVa7H
3EbkoeIwN/tCyPUfAQyYWcVqF9sz7U3Kj7mz3Blar6lZm6GSYo5/20OzS/usR8Er
AXnNUGRvPlQMDHFilHBNNhyPfHOgi2hrBhkxCOLNcSv6XXYS7yH+BVbopp78U/5x
nF7qDHEGO9l7a1cBtFC9M85uwSj7wkZH3n3SqVCFDCoWh21+hCfpLnOW+1l8DcC3
PrRXVspbdXZHtD7pTigXMEugQxsxVeBFbbAKxrxZ4Q7cS0ZyN+pta6F59QJ/zosR
i/xFYLBzvyphMmvl6AP9VgiSZxCQtIQoxNp2/snqFbUrnPoUwtY0nWymuCWMds9b
7BtMIqxvc3l3/VVJ+/Hh99gikOO0iGhAmMMpL4tV59F+8+bwb2XBh7lnlBN6d6PS
hwROEtYpX2nhtMKh+mkJ//MuwTjUUjzCZfhRKS2jebtA0S3ZE1GFYleuYglKCRAz
Z4xk4nC54zt41s2mHpfghv5j73aEYcQNqt7eO7+RZ7ukMhM62/egRWDQZ9cC+7pT
Wk2QtiJ6WaLdLw9JAbj/Qbkma+DDZU8xXJTcr4KuWn6pF43noCwX01gql1u+3oAx
r41ewSYKuwAMO83DBFEiI5qNBz3gDGYe2/SOGwp6YnqfVSbftksU4YutR+Pyxd1H
mQUR2AYV610Qmoz9whG+HbVUIHR9NBy1xClndx2rr42ahwqCCIRDSwhk6HdP+sxL
oNIqbVvOW2+xmo2HTjBrC+mfQICGqO8mGKxgnEJtOLfxxLk7EKVeKHms9wYUp6TB
5qLP1nQB9erZoYPKhCNloNB/yDYcti/wQJJZa1H2jxWxV6uXiRy9fyve/4YaOKyJ
TQWlY8ny0N+vykF6dUWkZ6IHe10Pmk0HWisxeEL+HlAr2kWhG6ca3OWM9QUizWA+
5HOMVBoxEuXagIe8acbMKyisbKSkVG5zyHuuzq56rahzEzVnh/AHxiGEbiX3Dm15
47p6YStAigJe0QFVcICOm/KYAh4oFmKQnY0tZT0LKhrLSjIY22f7Uwd0DrjpfGDk
CdnFEb8TR6Itxe7CrGICdqjCDGkIsfO/8ovIj6HnVNw2H6ZYNYYYkz3ueazhlD4M
X+YfiUUxask4kZiBM1Q2cGEAI59eQeMyZBAlSzH1fBxEoBraUtFivPQzDgQhYhl6
dX9QMk08A0zdp/fTgxh15mjqi/OqRy6qugmjpaUNoZ/aMbc9LqWp+J2rDRW7w6o8
/pbiGE1rQnHpjbtypRppaev/IbW3jyE8m3dRF2dtidqJnmNHsQEz3ih5/s9DPemn
b6Y2NnJSd3di45daBfSGa8+iebRDO0HY3saOqKjmTOl98sQoiFEe8/zpMhSpxP1n
/HY4FjyBDpPeTaegmdi2N5x4ivhas+y+0BTwanHlb0Rbb8ltUrJoGh/Qlw8j7ELD
kCbK58AP9fONi8CuSOdaqyRyRlWb6UV3txvk+z+rrIB4gycFRiGI2qVDaLB9loXy
gaj3jTnHeTzt99zog2tcG03tH+0OC9z0PqZOf6vAeMl6XVxaMgQZXy0jfG14Dk3m
+imEEDxLSaJ6j6TjxwiIgTvjxvbe1uOS3H5SYPvI97gFv4iuRcLIqpEYv73a14GQ
8raxt1PcLmzqpvqyqwi8WuvTM/KrTA9Ag2RlLY70jd8ugrhFiGanWQXIH0sRu+BP
8HczWwp8CzArN/aHNKTmCtdzKmeX5kXDgXbSWfW1yZEPkf5dUq2zGGn8f7ufj/Gv
g5U6lI/jKJdjsZ+1puwXBFhm31LryKa1eoKHTnr52f7U5YNtasv57YvndC4fh1gR
A/MWCft0G32/zSasDIHy8m3895dlOF88qej44ziBqSZ+q3Ca6MBoAyAflQmFfU7J
+FG20908Rxiy3jR6+iG+iuK8ezn92mDiUhM7+vkiS/16jTChsDMXb/snd21Qix56
FQosMe1ygHSjNmkw0QF8sEmKrTQS3Z8YFTDiXksshQKGJh/lLBF1QGEg4MgNNNV3
gUcdmO+rvKd9qGv1NXbER+f9Hb30Z71R+QYUmhkzlZNTguayEqfSgxshXJ8eL2XV
4fnrIHngvvpoS4PK2S8HxQ92gGIGqEFjmJg9AmWlnKW+acw9gXGqXuZI3rKLvvvF
ghpRiRut1iWLd327Zx2klVU5dQKgAIL0zWvCRllo1VQWKnvLlCxHgInCGhU/2r2X
0+mDbYLCqHauHMB7NoSU4sKcOs1NQPJPEb5ypTCI5h9fmPbHRHZzrmwMiRP+/hIn
+ArhaqanfhEkRI841V2R4NcZxHzBbb+fI6QrJOctl6sPK5uvthUmOuyTrMhgtCyI
PZ4I/8n5/qXnb+1xCE70ZMk74tNB5ELoiNMDRsiRzo5YJrpWzupuh0n2E27L0Fqi
RbqGnUOnoWMSSka/NOANeQstcDH+USW9lncFOnB4CNqYy9p874AkrE4A36P9rM0D
IS9HgqhsL2BmhZM67d2pjdxvxWtPkPrlc1QwRk2E7FADgA9O6DzHTOZttw4aeIdU
T+W2LJ+cwu4zS0vYJtjGSQFhJ0w5rkBuBQ3DMDwWMReUnOD3sTzRBbN5IUT3fofa
07gCLkOMsrC31gawDPY/g+QGSaUX66++zUCcoDPfLuHUo0z7URiojfCRNw3QVhgb
Nje1vSiBBdvL2V2GaH1+U6PziEtiCjxvo3scZUOcakqVQ5dPNp+f3OYoUiSg3kjz
NMDoGS+aVrOWMNOJwwwH/sYr7WSDgDqivmC7fVy6JrqSb3beL5AF2lNO4ZyH+txo
PM+oDVFK1qbNuBQaP/4p7axG1ETZSj/UAPb+bAmHKektxMzC+fcWnmMoPwhmXmc3
rzDFJGRHRUHmrNFAWY6hLTDRe/mpblKmHLjgWJiCbHQfSzqb28v8K3YKD9TnMnEz
iPnoMiHG1sBsVct6as82ULIPj8c2aR1v4mBB3eLPXTOfBjj7iWEVdcemkS0X8Nt8
vpuDRJltPUqNF+O2CjhKtnqMtGQTRIXw7z8JBWxZgdPXJ5gGrr756lBHgEolkWCo
S9Ku2gXiaZBi/tAv3YNYyKsTe+TOprB9WKN/7Q4df5xjo9D12u5YY6P3hqprIjhf
MKnDseMXwIsP2LahOlkH5pds6ERFn3TQ7n6o0pkgvepOqRxDZYEYLimmaNtnbKzB
e7kSdlAj4M6c5HD6j3CbdQ2V2ujQD0Wp/1YTTU1mr8d2rYIh/Sy5HHJq184IjfC1
a+SIZ0mGwvCofGq9rveDfcQ4nXzPlg1Y8Tn5c3hAVrUHu0tr0Qnt47EzPeYEJyBF
TII3cvLHd7gt8uNXcUgI1WVcbNwLSUqEOsOmQL+CAVk1D2gWl8Lk1fBY/EQyLYsa
28XoewZ2uatbiVIJDzDFh97Qeu0kqQo82ViMrwDfBnZK5qIcJ26Fe+/inqW5Teaa
sWCh6ZNvpdYMfeveNtBsTQ4tLRXdP+nTV4n9+q/QwOd/B/WbaotLkadjbwSJEwT3
o31qJBQP3o6feE4bnhv9kMoLg1bEUDwCceB9AmsvgywP3dqVKa78l8+e39fPWAMS
5fmBsGkbAQcY0mE+XAhshgozIpEAxKEu7wDr5at8geAEZspx4V+FD16S0rUmTI0b
4ZUfEF5V0J64yt252SiEaw96dKdihTh2D1WmATjqcGt/EpOrlR9Cuv43VJZ4r7Wv
wqEdppw8+c6omQiRdqKyBHhzl+k81spAzIghoLbbg9rHBKQUPO+bMcnonjFsh0Vz
5qO9cnCkC7zAiNBEmwqHgkpnc9lBlEUiioFkrwj9faY17nmv4twSVlTveOFsXSII
7sJreO33mWnHs8Po3XBgCbwlJBoMNGAgGt/pdHnFNRoJ/TeqPrkEvRyDI0oONWY+
WOn4EnBZhezrrGQVmyixtOGN+L53SPVJMpQvW9P3afMnVTCUt8+WQg0E/t5gd3H6
Qye3IEhgAdw+EyQQsy0i/PZFqWdxUiKRDmxND/Hnf1gP3WuKcUB0WMxsG9HkaKy4
pecXhWxniAHqcuNiG2INBxr4DsyIksniz+NlgItTnWRkra3MLVDhIIvNwh+bIPNE
VGF6+4KyBOKeE6vcBmte1LpO5jJozGQzBCf6p5zqd1ycEMqyhr2X2XW3yrEY46EB
hohJPJQiJg5oFy5oOQqosiUkcrDSII5vSsZmJsMdDrbLvJPPtpDMIbEG27jIo8eX
q1scQwr58wtEjy2h2YAWDW7mb6udDWQX568sF2Bi4W2hr+79LeYpUsgxK5w94QQx
ywlYaVLJMUVL9yZME2g9Q5UBPaCx4+On0wO7OlY1503nItAuJRinCrm64fTTmEXT
jAhI01azTRTJugUlUGJ6B/tShIEA1bOCBixQbbd5jQBd51YdC5xgiSp8I2rK1yeb
tFwLqm3HPo8uteaz6DmoeGdViqFhXY5dPGMQxkOyt54rNFc4Sh3hVC0UYFd8rP4Z
LQxB5VBcgz2qDJV0Zowbg3RMy+/DjxtExG00TLkZ9EDWwSnYb2bvy7j6dAS84hBZ
ZsfRzHgt3v3S3nNaSsydRsDN4NHTYye0aajTIYFeDSjpQIXgOs00D1J+jddJ57oW
hvAw8nkxnk33sarDpQNQskHuhvBfhP3Q2dexXYs3n4sb8f3r8XGmdYVtRk3aiG0v
jnLG+yvrl8XC3n+b7i5eqcQO4vGlhcOBzo920QUkmZZUAK+BzVOXDsMFvJBLs5Dp
GWajllPZjxVu/KMtx+adT7gb6ksf6u1GQJ4PmhEwLlNJoNzz96RlzcqTu4HHef0k
13axI19Ei9ajVrY5j1IdIIM5xi0dAcBwHc1P0F2BjT5IWcnESal4de8l1Go4fa8G
k3lEHmWbqj7S3jyQ6deDwh+hD61YZqRHIUeYYFaagGqhXfpLGoEeNEf20UexJcko
o/ljYOn+sNRjoPXFI79/bsLw0LFTmCjABhA4PilNbRE/jClDXWZzoy2I9vxSrA1y
GNHVdGCEPzu1/Ux99b6cEEBIMCuJUasa/HBj0mPpEIDAiaefW+WFBLh8IOg8Q8dl
24TOfsb0wxFYwM2LLr9xdIWcT8/nEN0B5+9c7WG4uNJrrufABtCbj3YxJ3bBHoYo
wOhFVdy4yJgY5YP/o46DMfR/x7OwBwzgKZ7jtVYe7tVJsUgD/MpeVIHBfLQlKOyH
W2qhIm5z0Tf3GUvmo0BAGYGU+P1lNCnz3bBhBOt7V6JuVJhVD1xHWKJvCAd/7eza
ABcaz3QmjHKprxGdN3OmNoGyq0YPTCPw1te2WMB13ayuNMLAZ+WEdRXvg2tPR7XZ
0zRAP2JHBIYWpRtwF5PQH5M4zAWLbcCQcyUZLePZjY0zWs3N4dIh3nUnesUtrhc1
SB+QCNuyJoGkFShgnFP4eoLhChvPGIT3+m6Qvhz8dLajyLlt3aECxRVes3Yn+z2a
ICCBdiNnyznrS4pJPV0Ji4cmGPRtNPOnf0/u/SZGwCcFv1fBEUA9qfPYtoq6J/ay
XDdbf10wge8oAHKLgO+B6sWkLVWCK1MgldemHZGFI3juYmer/ggrAlSaEQ/2NCgj
CAn22+7/kqNE3XM/KUS233BdCr4btOU2tXHKCyNS3gDi5QfJssnpL04TmokhNRue
YTk+FB0b29/aOToOAIJjY5ICb+dYvxg1X4jxAed1IGmey1J7SNaZ31Kg5aK89GN5
uusLd4fLeXSriKrFlaGNN61YY8EqnXg8JqDt4REd5sREl+1s1pVpod+QTKdQ0dKS
hYPOwRLXGaV4AUNt+/BLZcPPWRjidxZGxdxSycnHxu8R1iOWGhZ58EZnWsVyJYN4
DQnhneEJr93kfwsNld0aYY1rev9MqBpIeH6v4AtAsp/o+OGu3KwMXcMxmWsW781J
OaNmtFY1+qHc6w/11YtyqDRl8QT8aWGi5qd0zo/liyyh3LoeOXrypN+TzXJhwdlY
J5WE3oD0FzWB/jngel6o7fgCeNNA+xvmo/gJuNvVKNa8OLxAbQgotvF/hslYZo1M
QA8Z2VS4EvvmAOyn+C1ESc6fhg/fi++rK/dcBo8gaq9nTvZaYCbHkegtprMXb0Fh
+Ag8OIN7iVLhu3dOcw4BREDz5Irs2THSoTCJwKDRHOZsFr7lxOdGNw5UTdZbWShc
neuVD3pdsSjby3Je3pr9iaSXLrh9XsKLf5orML9EE999FLaAc8eZPI7P6lXbxX+4
Bg1/jzLHddQsrWbWesMXgcKJq4CLf6E15ZmVpClTZbXxTMcbKoBkZL4aJIDxFeAz
x6lcS6Kc8UNUCxI5WhJqNwiSN1ctVLhusMq9Kuzx6IgLJ5CMUBmETru9l+2HH4eR
MamqMsO3t92XLJYXIj6+nHLeix62QcFksssOtH5ler7xtyu1H8wUTuZ5r5iv1e4b
SNvZhHNibcIkirGFI9eJKWU3zyknutHxZGMBQnn5zffO18CfdUR2iQXLMtz6XzR4
/IEEkrHhJGrPp1UrfiqVSt4JQLvt3POaGRxdNwo95N2eHIFDDdmxvtoWyxolLeEt
fV7zSTcdz80W+gnia8CVebSvR4NiqsQTZy/rfW6P8l6hFomiMs9IFcK5ljJb02yZ
U6vUic7H2INPDbEX5KbSSwKcM4E0AJJ7qlrDHhZ47bg78+05qlvhMPilSWuV8+92
1YTyA5SpzcL8C0mnunCwQu6u8hjz4CwGg88Wrt2jrF8/YH7W459TOSbwEsGlp4O+
t87qCmG0YRxc8gPR0LI1Gee2+NCeJQ0JyU/WwdllniXOlBewP2lSMUyb6ITVrxep
jAzlWKRMAtp1XWEivdVa+XIJxtpJjkxE5Ym4Tuylt2yjxzrnXC6jeWqbvRVNR2QC
2AOHr3d5Sg1fX6WAvcM75d9t7r5APghGXxSGiYi+r7e16UxofoJOS+xhYhMzs2EY
0NPdqAmqljvBEA03LR8mLts47AozRot7Qe5Nc/X4ZlM919rbsKlH9+uEkB86keIC
ginOpyyiszEMKkltbY4wJheUd2gJJdP2JD3C+IqZytLjHibmdYZNunOqvDeIOt6c
0fGymBS64f5Kd0i2sYUTxD6DqWunWf4OgP301fy++PuXAH+d3caklnqr7MQuGSd3
2BuWoQLtQAXeN72DRTHxLHPCXIIAc9bJCZ958AlfjfTb85mij7PH62/IidGr6QQR
U0OFXc18IUyppnMy1mFZvHUp9qzc22h6hS3++Y2RvL+KhevE4c9JTpoBxTJ92g9r
C9o9kD2hykFstmdGLDp3FIUcD98hrzUKQtsp09y2kdgG/od/aprlRLmZLsdIx27M
5Bi9NvDmb26KwI40+su3Lcx5IYQT1NA3S8+TF+rNgnlIv2Q4eN73PuZeUQmQa1tw
mIiTYEF0HHw1bTccLJ6zH1rcevLCSDOde852N1aTk6jdg+lVIecMYzDg2CqbGVZ2
GlvqnyME4ERd5s0v2Q7hXFQjOzrDHajoSCSKO3uT3GTXTkSbZ7hRCKn+ROgW+NE2
TiZK4P2RNSyeuiuZz0aDxr2ZllRcqBAPgKaj2iJMCJGDSzsZGh9phx2Z2HNahyLM
d/tQQFSVF12t0Kr8yqFECl3trDUelNG7YfThVWPlyLV19VdZdGA+nNEDu5ZXVomg
xzI/wg9NPSrAz+FrPvEOWr2DgZk8x/KOhe6sHIOonF0kyfqpecuk5MAoMo6yVP/K
4GYpyZtw6gtn0/M1uihSwG29XHudvQYnvLTSijBgm0TkKrWuecN0fARQBOYK8PDt
cFAxrHQatb7Fz5MGeQhzLFQnIJ1b3KGij3qdjYO6oDkLjZ8TlsGI1Ae96TDdbdEo
ZuCbQ34MMGMu4c+YysuTQgx0jDeGzU8u0CeO7KyQKZTXghMbS/IumWX5Jqga4ORJ
8BRFWM22L3+uWFgPUwhqnEZ4/LUq/O7aXivsH7rwkXOVydQnJdvVnwMFTdXj1R3j
XgKYwAYlPoInHe1BetEbRrFF+tNgoeAL1ZJDpAHQVF01VQGJNbnB/Uw7ki2zXR7Y
gYjnzzKesG8f48C52o2nLWscOBETVbAW9g3qxkpntb38wakfhbqMpQIFwOrwEg11
0ku/5tYfMKHb1HKbt1ni7h+sYX3MDhIpEWn4rMxOXfQ5/BBeKIgX0rGrUamMmFN2
EOrm26/hydmpZ8PiSbHeP4gWuREfmRSW7HxghiYpbdtAt2mde0Z702ZFCiVItZvM
YAarxaLHUJXGLtXRgmhUWROvIVq5b0fUsc/yeuHT1EB9dUNdNcXdTW9Vl7pITgk3
E8AL0x3BZ+UEE8lJ5BwLkZHBjt2Ih8V9mcfvk3IR/yCYMLTmdTKnTnqK0n5mOIyc
+Hm5XxPM0cwvMbwqRlJ6gGkGV0U5ENus4OmSj5YVUrsldHK1jV87RcXQ+ds7M5zJ
Y6m2Vmx5g/u1ghoVKtSbYDT1Ho5WakOH1lzpOcFtvSJK33yRf/i2dg17w8dzo8sp
AoBgxob3uDnyWJHN6X6xoVp3+PHsC+HBx+BQvBzrWcL5wNMRXNdK4bM+sWBhB/6q
HlUy6fO1cAwexDhy+F+s3nfzo+zX8HxS2LtSCkIq9fLoyXh/oOmza4RAO17qZiux
BEHiDOzkrvggcxNpZmxcoZGWiYRyCKq1zdCNKs/FIHv9Z+YNzHovhQnoYOzAOUMA
WkzT1BNyZWtcijJgXxaORkAJzT55rorQrUqHzlniRdaNDnqe77FifXVAUKaAnTYd
km3o+6klL6O0/gwpKWW2mg20s67erQBrwsJzHFOJwoFZPhsLcwPYt/1v1q1R3OES
DHbTcllTy40K60maS9GOacqGlF+2A8tu1lsJ4TmqpVGNpMHn/fm9SP+ksM+hRhNh
c/6yUkaCsWX00xW34rgKs0T3q5Y6TlZI0w/f4ijS3mJ8An0K9qrW9byNVlHBPo1K
N5TniXqwyXpuYOTIZlOnt9HhzZfg5LZtScOOVEKcCko+U8j8yIWwxxFtjWrWCmJm
ZlIMJ3xsbImN6n/DQyByxf0nDdn+qD/N0gZ5OtA64FcMSlWhAa+/huwdV/FyqMTI
8be5uU85ve3dvtm1hs/QEgLWmeSahcEGMeU7rP+WZm5Tn203WybTouUhUFlGZyiF
uwWTEWy9eVfo24v8tmbE9T1muOOMMp9fDdpCJpKukV+olhMfX+o3LaAIWQPEPNy3
+r9MDF79RVL0mewRGNmGxDM23kWgjDl1QRY0CF95ou9zsHy9H17qSiTca5qOJbMH
M3vSvREAdRCms4csDRqCtvG+kAmVuhafui86DccVGN/CFEmVFdD+YLGM1gVwrQPf
gAfEkkV9yzES0PlUNBZ9O/s3mfjdRvCwAShiwZwnCzn4HNx+ekyTJ1dCjwA6kRXY
lbwiUQBPQ5+wuUh1p7EoNBaUgSxV6SG7b1b3l/qhA0fHiSEWi2ZPAh77YuzJJQ1V
9pKqXsrvGCHZTOASly33FvrJcDqPFGYXQGexgzdbs2FKw7waExzYgIAbqURFA+8K
p1Yn8QXFG7s9WOCbLmhS+369mMAP6kbKRWgeAfcZM17dyajoQkzmCDGT2M7X1ADE
X9TENSkMDNMmhCAYRUnSmGwLPgcg8gaagVP1ZGpaz/BXeLzWXnNp+efNu6XC18zs
0UK98u2VsY15QrzwaKmuZeIYwzXb+ymPFJ3vmX0UJzEbOXtqYJNg26oSmTCU8RLm
SxBwru/KUI9btX+vG2Z3KfLDUtp8kWuIBZaXc7Ras4vOtQv/WFJh/XiXjCYEwxcz
VHQMGsiJqogceIQWig2g8Urvl7ASBIc2sRVKtMJiUayUJ4VU0ASArYdvKOWYSSak
yySuEGHdn0eBNfTkw56glrgnvLSk7IUJPc3YzbgznY3euR5W5izd2GnjJ3Xgb/Pl
2xlh1a3Ct9049AgjJwOHt+s5mASy80uYYTJad8zXApoWeVMiKPpsBE10HCsgsJEB
I/KZVr4keAf/8gtUZdsgfWrksirm/+Tdj5kQqwDO9QGobJphxP9uP8MWVMDWylZK
Lo0s8Rpo2zkUaL7YL+TnnqIGVGYljl584wZSWTFO2TzCktQJhY/LlenhR2sBxQe4
iRZFTrL2cBLr2VibD0i0UT2LnNDP4z7TXC/PcC28r+jL79++zUNNxiBsyhuHaNtz
6LUlpJ546xVoQmPa8/TEiM9EZ4Bp4eVFo8km8nHNhZQtdvISF6zf8Gb7Ypciwyve
8I1J3vpXz2xMGRY0MEj3H4B7LugkFUSPDimG/lOLvEJiiSkeWoimrPJgKITykODL
3ZaR17QYJaYPnlwbXfWtd5sfQLE6r7oIp2jWlBf4K7TLcg0MGJvgq45MRnJUcWsN
v6Rxuy6Wv6apKOymsS5In/lwlcHP4+4PrRQgdxRdxEW41moDAUkagkmoL9lwT/Bw
CrFccx+up+zj/tzIlhWtSNO32kuU4P8fNHVTbWlJuelGsjF6t3c3Av+/Pn8BZ+rO
spnhzMaCFlG3C9ZvoXFlS5HoZ7LaGhU4IFQMBAHEAuhkS/BWq+MlGU2/4au1zPLJ
kHK2qnR/Wbg+zIr4n3OdFiravVyZJnzMTSiCIl1RNJRP7KY+xbCyPk+ovCoGvR7U
1TZScRl1PqEUFnlEYkfyHMPyiGoCcxmFlr0JS6s9yfUUVl5t+rnZGT50u100QLuk
tQOXCjY4A5pQVk2PVgT5MCEwD6XaEZxSXuS+ZY8S+VHj/4vbXevbhT8A/yEtGEwB
AJCr+cpfX5BaxSLg1ELGy885/V+PNjkCORGft34OgdDittovB5DVwX4lioJug+8B
V7yMyJm4j1uC84K4nG6Ip9iJCtvJPxrfZrsb8TcF86jqxQSTiRqjiB69mjlvz6mz
HAu/9hUFrErP636D88U1wCXwOP7AseTlqbPId9H8By/VNpLeA0lRcXi6d0SABROX
uxYdnMADDnqCy218G61pH9gFKGGR4jZtRC0zpLCINjeOpBT47VYWYGBNOOo37esn
9lKDoamartvU2bD6L1RiM9/rg86ZxmkItZ6UigKGBbUfb8Sn9GErFlBGiyBkmyzt
rWGI5yU1ToPxZtTXADuZ/YNeKPf+j9+JFp5V2Z1aMidjcxMWmTmWMqjhP4DbSEF4
OP91rRBzyJpfQFKQvqsjcAyHqLvIMamS3TradcUtJO3wnXpfAqln5a05BETNCwqB
xMIBhaoEjvqc86FmVoJa2tV/jMEPvvq4BtRBhhbE2UfLK67A+VxiOyZ+c5ZXFSno
46Agq4e6maM3sZUHqDSUbJ9x2JZLndSPpJ0Pve2ri4QWmWzJPthryAiuMWyMA+Yx
rK6xerLJ+cbDDCYSRvDK4SNiFX/x/CKeEewyz4eg/lUyomt9a6a+ZuEie0RHiFSf
w13yln1tj8cV1RG4PL21K9KE68AT9bFQnuJAzAtCxmdYfeKnJ5R+DkI7Q0dAQn3x
1phGqPNdWHSdh+e1/NJljq1PuS0GJ8xt96GMLKCX1X7Aaq2SiCVDYHOv37enm5Wd
5c3ftbbHyje7RJLwB2qrd0kIGHKwqrbu4zKqwXg01ZwQH5ushMYUVi1zTWZeDY+A
7yol+cOVesb8JUU494y2nMgHdAP5b+SEHxth/xx5SdhjqInV8ibeaDfT5Wj0VVGJ
L1hDgl+tFbwNWUpYn2Ven8sbp1d0eg2N5g1DLVzmfbsIdgpx+k7WzNOjQjWSYq8V
qppf4CLhQK2wBRA3jOwiAY14OWL1kOtMxn5CKi32sPqCDGtu/7hkZXcQRpjR9SAd
BTAtRCCU+BKEJZQ9yWc9324eILOcFAQbivH6BStlZwMMoVcdhTRSbTj/xbjo51fU
kdPWjWTKpwQu7UHrnPzJ92qCjKWQytvmli0T/S9kLgr66+u7owK8v9KskeWHRxHW
IerA+m2maUBI7oprGiKOE8M6PTxMntzyF6OshWv++GbudvBbMwcUIvjcBiLLHoqq
f4LjdsSuvwdYFRdnqWcmYLXzx1LpFfvnd3MotqwTGywKnkSlLDp6Bo4wtcAJfeGG
ye/k9sVFYZk7+/dsZql5dHxX3v+HsjogiCYZZl3gb/lEXDJn/Ei0ZuHxjy9M9mQE
pY0ToZb81jFsIWf4sL6CWV+0+/0Z+dr2VAi2vX9w1aZ51/shB5yudesGZhygUkQC
wrm+hz9zAX6+CSz6DlvG6xlfsaems7Y8ucSQdZslrEuUXx63Cy3sMH7Iupa3RpAZ
60ozYSz/G4N6jkx//XLab5VZIY69WzpcfesHZD+Jh57YDArDmowAlddJBqazvfue
ry7nELHkdayWNbS7f7p/6h+dBZOK5nCVfLCbMTZ10wLN0jjQNYWuMaRPG1SHx+eR
pL/9T1fw4yl/2Fy/Jp41ZqA+AbVEMv4wDy9ZRWihW3SaLv3Njmmw6ZYOWojhDCPx
A+/T/BImPTf49EB3gfXQuRvB27cJKeN52BEpiPIak8MGzWimxYCdytcEpkjbOaNt
ZqMQ/MrofZNVGh2g4drWDfYleMKwVkdc+eOrvQO1ZXxGSl+Ydxz+TjPe428IAsoK
PVQTUGs39ZcnYPEYhWu9nN1M3qTPYfJzSpGF66RIw0b7D514EWTwdKioVZE2tVtT
VJPz9W/FRr5N89rhTuGtG+EP/WHQPByzHqI1MiPayNAuHwVggWtbVRoGbyJTLgNY
DFBwy0W76H3C5jFhCndAQnfIndcgZRXK2TB86beXejJRzdSyaWoVZvk8w4qLcygd
y8UTC2pngKPt9zeaVQDg/A4+pJzHDCoIHVLB55zydRGBCVy4TkZ4zDg6j/4LkeoI
+d7lno2FV8qOmsvxxijQdtcApANGJ+f/8OrG3zRSpy+IeXE+voUOhvqNrxmaZ0m9
XY6qAZTgu/i0Bc6mDJwcU6NMNDf2bbBUCwsmYysegiSboTdZIB5MJENwFC8a2LxX
7tiDIFeS5Q5KmAdo3wuYDYcf5QCw2jS3T5eR3C+AiucDcsjKQt8BJYgZsJV851gk
LdRkaUaik1B56Dxlo5z8AAUJbghO+pR0Snk1UcABKcm4krncS2XWsR9PFcItZDpC
K3qU+N6SJW1JLmAFEJtt3QRTLtvBRmgqa6bEbrCH0S+7knAWcmtUnzlBhVvh6BNV
efkfBxIvXkyxtqhVKYAI1GbmZc04O2bZ1o/6Td0dywHp7rv/at0YMp52a2YE3a/6
3FarJ3l4Zvr/wiVd9H1w2+R2pt8sX8X0oQZiGT7MSYLW++VYCcDxEtHJlaALCeNV
n2obbnpHVfnJD2s0eXmQ2uJ60xce+11uPsiv3v/LPl/Kf8Kc5EIckh1inytlyLNi
FbmuNa1jrXiiG9pYnWunm4qRWU6yUqV1DvtqeaM9WFRUaiQvUcopG70ASmEoyPSD
bVTQMgHjB4RX9o3h5vrwnhekvlsrv1K1wfoIjtaK01ouM9I75kzUz4lqJNhFhNh4
uCdmqiskRjvVrhP71GuWI6gk+0OmCRwISNfRA+XgucWzVDy/SIXUus2FBKMXgIm/
FTVrptfRPVSnSJqmVs7UzP0LP7dbVY8NChxkwIVAswTRiJWLTXZiwUavibcPvbFf
YYG753ukYIQVK9qG9Ih0uybG+nM4nGY/0aYmxNHaS5yq28b9Dr7QWgSfuzUzinhx
4rN+fo4BwHYfqjNzdir+jfuChU90CrKsWHWo2rQ8RJT3f+A2XorJ0FJhMYW7KzsV
3asO8FeIHafwu2BEuXswDycVVqmZa73MEnY94/CQmgYirSNwlQk+FsfGcQ+2Gjt/
TRrpnMfjcJxFC2A4VLBjeIJZbwfAvKtTUjTLERpXZ+roy2DKPlN87hVRZAJ7ZPc0
eBv6aKtzlOo3ZyKhGGxu5q+6sHCcJMsz2ZcqNIFYW0QJEXzdcA08LZz04lRkcG2J
KYWJZNZ0a9UWadm4J+xb06RRPDL7ev5WRyxUqGpiZKbZUEFj1L55XulhU9o9EOX5
AZmrMPFzAfq8WUy5jMM1EpvJBJFAWN9RnNLwoqYo/UEDffClRcJxCaItUjDEifqc
+Pa7mRmGEEgEolS/AjClhYoyua+FPRZTGpvGkbh6uYdGEpy4Yv+CdfeQvUPHITrM
n4Fiaumq+/RHU4tm+7noy+731zVJM6mfwwVeK6DzNFJR3LaBqn098GqgWUAsnQMV
nAC2tAFRVe1tbPDeoPu5KVTj8wjbzntIVyCx1Z8ubhVn4Gm7/52B544FnzCK1Zj8
sATCkmUc5ns9mhQiTb4O6aNE3pmxOVsyEctMtOpDga+AnBGnKH4EKvLniuANdSKf
ti62syhunMW1DvN77gUOf2RRswRTNuBh8uMuSwmv15lEr+/tdi2YOdRFWt+6ufH+
6Uw9N/webdlb7rLEpgDQ1cO6LTebvSefOrsTooH7lY2wz3REv8D9e6x7KnMFuZlT
lthR0pwUY1yQm2eXh9Jmkh9hMaZi9YW6DkbLO6Xi9Sl7va+pG2aq8Heoab4hH5iB
HTtQOWxr/9IoFEsWglvBRBu8NjkwjmyhA7bE/r/t9XCEFpt1NSv31tFarRRRs7Ik
EYKX6iOvy/j+k+uUSUHjgDQHiHMQVhVCJ2HQFSdIynr6kD4p03eqUkfGANFUkUR7
M+/svvKscQdam9W2H+YtkxsVzxFTabUHzo/bT24qFqD+yZ3qTFPY0NLcbnlC65dJ
W3Q7JVwrdkga4950lrDnD4LdpbR0Ms64VQ9IoNqdn+od7Eh7i3D/oo0CgwV7TnYS
w2WWHwSTWzRF8AfqlLPpLn9XF/6zdPtVzRAgEpTPyIHsOlQgVbM2aVAiHtF/sWE/
UUDSbz6Ymc7Fgn180lCKEP+dyEr0uFsTgxLEn+s3Z1BrCpUdCbkr0bGL615RKkA+
et5ClFm9nuV1DBN6s18znnw3g83BFcOM/vHBIaP7vEdx03eu3iBWyP7+th1I+vFE
8nf6ltwB52ZFNc9NWgl68wM1AdadHZ51pgCpws8nYaIrWOjf5gfewPlvhqdwtuyp
ffFfObUmpwFGkzGXGZ6z3WvBDS7UEB2TOvLIimhgaKOuSfBV6c1Rka7xHcrDiPvI
g6acmgB7UnbgrMw6ljqZk7UmqVkL4cRrDUjv24Gwa973eqxJa4zHVoxe9yw9B/bh
XbtUlCtkYjtfCZaBsJxzunE+PZGx5Vr4xoId88RfJfDjlUHOpD5YvqoDjmPv9Eta
jDiSdGfKmTr19yLvmNvjJqK3mb/fsLaG/A6kyTeGRdlfgHnUhQILau2cC+lRz7ye
p0Z6Gw+ieAqv1qlsWhfs/r4R6KcfPO7JGlAekhPTGvGA23A8u3yDDI4FMtYqqfg+
VMtK+yPNWNNPukD+mdTT5JkLKpo8BpNxkepGx3wwjDm0BqSqPtzz+E6m87kn2VWP
krlY1suY08nqfRw6dupahDuA6VgqSGR06pIkEluzujNYRm5M9+FtuBMACFXWFd9v
S7rYSe+Sv5t7wXu4ABvjs0YjhScWX3S/3KTohXNynPxqirIiIfAY5LYKpIoFZuUa
v2ZRFwSHM84yZVHh53p0RZawvLeSM4+A66Yab9VbNz4K9bvlwRrqznqte49zadY6
Pv8NSOYZHTgi8+LRPR4osCgWy5h68zl1jvq+G5ylOaffiQIgz/0UNwUOubiDOvw+
strWtXByxEEQTccXuhh8QgcHId8UZU7X7mXqvSUygWl53bZRbn50lrbS9et3ZFPP
cEI7Gobo8LzVHwnQHHaBDFpYdDGdQB7v55TYZgdPnYL/JI7DBVeBeF0SJLqu8DXx
20SKejkexwPKbr7vEKg/86FB8ZsW15HbRdwqWfMBijdtz6fjRujkrGbKQNqT+c+G
eI/TMD/wX+zeOTIhL2WQHKobcUr13BqrAZTaSkq+DvWTjszXFpcs9ftX86SBxLpz
nPdU8pyUN1Whi7xi0qBMOEtLO8DuqXSRC4JhSgNYvrfd0H/BbyjAF6b7Ikwmz97c
pEJXb9ttKp/STbGnMZ27fH7vxrKcNSf0RLnZllg5eyvb3hjP5Ds1p5TKq1rMTj/I
8ILD4Yp0Cv/KSbMgWgNSmDdqyoxPeCMYmU2RwfV94XrWVqznaaAyhqffB1fQ3Gxn
/mxBuEqOaGp9Iwgt39PxqLm44H5v2ToNp+kC1dkluDEMz0b59PtsR6OG9cqBjmRz
d7fEJGwTFJC3HDyNUkqTpvroKCNnCYREvw5MUWhWaRLQ8BhpRGAQZOX+wvVTI4SI
BX8cD4OeUNPFgXncYZL8cVQ59HYa3ke5kiAL1P1jPwsGKp2fc4KlF/e8cjtn7HI+
TuYZdHpfwEr7Of5NpuHP8mEfG5+wJBOjnJ2FHJiGYBggBTvMmLf2RbwBhjlinZVc
l4HSCMbVDEVsI32rfzxvj93U8H54mvdKaVI1p831lsDXm7otYf2l/k6yaBhD6+KN
51tlpncqee+vVMnXHMdcNslz+J1Ke2LtC2LwNAtK3drqRlt/cP5/iZl/+24lGCmV
yrXFkAvlN0/FrbEyXaYWfPhfNst3bHldU3y92hxQqSSNZD93DXQVRdrxCwR5j8gC
eFXO2vA8zu2m6kH/RLSiTA41O7nQ/09UIDLwzl8Sau/anFW3h1yFO0ddZea1dIPN
NTVdU4qz64UA5x5DlQYganxwG/uWxbwm/LGSyoBTkh5ChMuT0YdmSr0SFeI9uN8u
SuS5K/19FWy3yxyIDPcp6xnnALrZsznZjYwEA30bNQPevuSb2+qDvgWf4wGnQd2x
km1+MqHuNFBqUHenZvO7rH9FvKR8Z9pXEPeqv2/JF3vZYngi6TY5hQJfT/VDuZXQ
W1LmBDE7QTWkWyZENAMxPXFQbu9TMTb99SLadqv5nE99U1e56w+esEtrvref+4KA
+iNka0tjIPWISAO7Rz5JUimwJBp/j/AKdfdGLG/Y1XJCQGfxE0q5/mU7JfYn95+j
HSTLUgUZG01/kwlghphIWAfApQVN+8Aq6Gyh156rQzY0Duum4hVZCLomGOxYWv2u
9j0ax0MdHG4EaJ41nUPjyJfYZE6dtHg2H+BSqKXtqXfga0MWyWbSR0ZcuY1a7x3D
HGI9seUmkawCivjfMjz08djHd94hynkCaxh09dSALOZ5PIVpoxqv4/GVZFZgJl0s
+VxcDSRPedhB7+E23ElNKTRVFlFeMg6k6QIRRq18k+LL+/2fRyhsfRz/U8yNickW
yUF0O/I/XqAHiT5SgHtME8DM9pGhLxBliIHQTQ+EpxS8hwBk+uZAnO65mHz8Oirt
GNPfz4sFqvf2ydihA1rQIu9TyD7oDZzaGToBZOQxHmJmRXwK/01H4Q5dDKKXEKjF
i4DUw0YhqyITIvrxNAIP3/oNS6JccgQrttGR9W3rJJwEaPYQqKmyihakVSt6/gkI
umvRD75GbdecZjI9d1vuTrbkVW004Yckgh85dfIAHrbnWfMtiI/3CdH4srR+lZvg
iyO/X9uV5VM5jaqsjjhDyllj5YOysh5ebB2XJvIgMygam3yTFrQVK9YzF4oMxl93
zPaeCFgVG8PgS1xL5ussxXvSJvR4vH64m4iH1WBdSiH/B8a+4HO0vKvz2q+B+etH
7gb/zrPQt+stuHCLJZrfTrXnVrCZZZXIO0P84Nt3Mw2ZB5x1KEYJ4EkLqms5hEMP
XZktq5rpARBhHZJRR4m2DGS8g2TaxPSHSH5miLGK1X4hKYdZkxs6YgsUvDqdJVw1
5IZ9w2FmOswLHmTzHNl7XhBFfTh6XAl6kv+ancR/auMEsAjSvCAeqo7XuX0fNO8C
4O+LdTx8586/n/hAGuqkDPM/UiVBAcWqMS/ylkuAO52FPzUOlCtzhpfIxt5B7SEE
JI8SD2unhODf2ln3Fy5pg5SdrLmqW95PDFPIO7RV4TA1yLm/YmVNiUwI4q5arKVu
JsxpzZp6nWo1/1ZMCmZ1b5xtMezr7bcS3VLZFEZP74h9faoilmpYURKDCd0VJGh3
HItsrlJiknLnoVHmwMku6hBqEQMXV4HOfAbjHh/jZpsQy7JiSCT0mW2UdZOX5s3o
dc1xtsm34XDBkvuty5DEV7ibyWu9zUmzH/Xs1gZXvVUA3054avfHz1SzEumxYLn4
Lx8FbAzLKcmqTfczY9iKLYNpzupr7BSu6TxhFyJ+5YKs+oE1wQDb9Mvpf7QsHh1G
BU7CEf3/Q94Fd1u5IzlUTZcSJKSI6IGduOn2FPVjaKWJPAN8KQpWWFSvYhp0NYuf
OGhJ/y+7ZxT8LXBiY3QLdi8tmEEvPV/FVhwKX1SAdbeIInb5Mxer1uFKXVhLbQfO
3KLWju4Vw9575ps86FgSa+zn79+yPtS0J2M1txOKuQlHwa0FA8h77IUg4Thz7/S/
azX6PDhbaJc+CvpUzo1a9EAIXoD+ayJRJE8SJPKosfi7Ph9k6RmFtFSvkJ3ISAyc
t5DwdkAt9o7KzWtmd/mJmezFJ+VFPfc4KJObzbBmRcXDilcEt2z7g75IX6LqEnzU
B33nv5XOnUUsA76SEXrqnDybzwocH6Ir7KTmVFEvVzw3GMeQYaFyYNwMfxBG7PeR
tN2+1zmkrwgHD/J+Ffs59s/QLVi4JAC6qYOGXo05+K+/cePnGsza62XaTEDDK8uR
DNzIKgYXli0pSD8rn0zihl7ClLHJA299pNnsjF8neykZYjRVrIeA4M/+AN0rmBjC
XFU8q0wdi2K/f69IPlX/6WuOzgWX9MJg8FCrWhb4SFvyiUYQpdlOZ20Z0QMyAJhe
JGXxaikjik0wHzYYYEeN31BlUkQfOrAKGEmP4H1IXpAN4rVILfF1aVuJaNuPMCYB
oJAanh25K5IvxzW/3plCVWBX7XTFkH5QeherLgLdgY5nuHT6vJeLSpbTN220d2MD
SnwmWqcDt402N4aLPImUyojYs2JvxkIdHnickhzE4q4biVNOZFHkTwiS8DYALKYt
Y4oQoqCmysHTZr8w8DPqsKcF2Or8IGMKc5k0ZiCHp3IADbcfEMzKgIWcjpce1/XH
waWU0a2VRw/7jpSKcZpOx/F5SnPXUC1uhZYHgCIpmEGq/hOZAtJjZfDUWG8+5xkG
Ofe+5LLkuqhCEcDreB+y8xyhDbZQLbAI3SWBev6wxGoZrN6s4NE1Sy2DqJ/qAFM3
xf1/AvcWaGX38eTWFpV1sZfYkIbVhsxNTNS93+1LS1+PtzceyXK+xOAivSGyaPZU
5P76aB1fzudaIJQGswPfCfRegnJUNKno2PIkgPM/OBrpJC4zHVqN37XzijJCO+Dc
0mucbHyTq6MnwsPyurSrCErqYgKI0SM5/Q8PWknkZIiQIurUDn7aikEZchYpHyB6
npZXm5FGqiGofLjkX4oaAlvIpr9YFa3HKydjupzs4MEaBxO3MI2ONfZyC7TUwjcQ
2mC/SRfwsSvNQRjWM1JKNvxJz0vdmcUT1sKstkQBs4YNoIjEtU78dk656XBZNYW6
t2yUDBFXzzj9sFt0wArJLweMz4nsUs3S2YacYdG1Q2iT8hRHwu7H1TZqg0En/Gzf
vny2OSpFOotqrfZAT60IwdzGA8eUAc0K0uOujm535dt1eEfj/AVvnF1Df0Am3FH+
zSutg0i4SB2vFuIm4hIZqKIi6yZCc+fFFJcAflT4HitOmcfLdBQeqnPq76VqxJ0W
asoF3BJYFbp1FIGbYS4kKa7CpsY1wLncDQjnoGIc6UydmMof4xp51PcPsL9uUt7g
6i1GAbI0qbtJUkp5Mr7Jwe46v2EJEGj3zlIFJKZpq0kPm7auOOrZmhQAc1VKxSqe
1qEsg/K177JgdIXZIxyG//tql+LwPUgDRR9ro0J9OLPrQN3SYOOju+HKqDRQqNdd
8/tzqjSC4WLzEuFNyz9C6G2Bu20WJX9lZXuQkOXATk8E5rwOvY04tBodDL9TQJqU
AaEefdgqTKLFlIusZmhGofej/pue3svpH6UzLrXGe0B/F1peIHlnOyyU0dpNWa2m
9aLCH2IqYOBvOK61Nm1run1MTpe2W/pF9qm5iZTJJB486N7aJZC6cOoaVTgVONBO
w5zhuNISerEbYM9Q1FACPw1vKCw0DlRlGaQc3114oLo0PseulTBFDU/cPYoB6JJf
QUGDm9d2TmgluaclqU30EHOU2Fk5H8Xogi7ZGXAaiFjdcG2Tebi/FQNlHwGr5urw
0Egl4belCcgCvY43EM8zMTE+mxyyv0gJduBwqhCLkD6uiLJweq5qS6jKyeypFQ1G
B+FqFr85ziw31vKzue4oBmJ1eUczKwiqjKu1zRwoug5QIOb7n5vUk1DhvPegkWdt
1eYEafRm7UpaUKzS4y6qDSLy/xotKab6SbLZwGSgsnWoDZjhMMS0X9II/xX0Pgw8
VPrsrqMXFcsUggZtzxRriKgTkPMnvwzBwGGjpHn5Y+lszsr6eOY9drfh4T5xHtVu
8NtW+l+Yv+F65u1VFerdC9mU/hDAZBNy09pmJgBwO9m3WYTSh0FTjLKQyz15vFfA
EnIvbSKZR2KLt1DZWNVanxC3UA/VRoMHZS1eh+0TpMAswSwcHt47xnepdO88mcR0
RnOSGo2bS8ct9TD921XWjZpYydtcOXRuJKUoZr+H/OY0mfvgBBe652E381ab9ezt
mEmmewYuIKsqXPIDCSG6uLL2pJ8z06v9H3Sjrdf7e2SGkG0SZpZ3jLurwf1VNaTE
oqXH1iKiwZvtpO16PJ2Z9YK7hwRA2yV9OSCES//WjtITB3KfoewgaYID5xhvv3c0
Yu8YbGwb9lmVtvprHL8j8cVaXSztyuWVLMOAgFwJE6Xk7Egi/qfXrpg1rdPVB9v6
J7I0FOCcVTGR4lUWefJYSs9lu+6ggWG0+nVbN7sUPvh9tH0fslTep+YbKrqKYX2Y
OGtdGrxtnwardDZ8IAMxQy7yqDmGTpHuSqXPD6eg0kFDuXDq3HJZJ71yzxT4lAEx
fkeZcLyFsRZdy/JHI0eK0e3h+guVJTwswhFAs8wu6KVr8dPiB6Do1qBAp6Fy5ohx
HzntrHoW0NwmAnjQPstCg6/zE0Xmr9xXz7i8OrYGY76mrIMCAKiqwikZSt8VDtWr
5D6/OzVVbybGNQtNmqbbQDnq5Oxc8izAgStC8558ISey5QEQ9KjU8L/xPd9zJoy/
ca8j3fGZ3cirPCuOIV5lTssYolOD87FSyL4MTAMWTGM8Qo9VAI6Vmteu/DmTfsSu
ZM3f2eO7njbEvVvQPFOWO0CtiM5Vn1VO9YluuFuHyLs9OlBg1xYsKd53OVPjvqfY
V4p84SbSAWK+IZcBdzFqOJJttlX0DGP10KKo+/27XZWlUicfL/VR8DB1LylIMl1T
zZYssMBMZteXlGIwYN+HjRaegTUcN1Mv0nMTj4/iOQ3yltrtcC8iTsrQ8UmQeSGt
22GQ7hXCIM+os1QN7g4DiCzbr6y0kNSQWnwlb2xoP94SH4ttp/dEW8kRvDZiJu2J
dzGWpeO53sfzySbw3e32LRRyEkFXVSo6kiJ0N+xoRkIfsdxx4DTqL3bwlNwVjAog
zICMMDw4MzR+AvvsT1dF0e33gFbQA4KRfYsIJesXY2c+3cv2roe5x5s991/GjB20
Rt3fECotQwhdb+HLRAz9lBEjwn3fXtV+DhYd3Hgiu/rjJFFC+9YuvtUeq4YXCczj
GykKuy4yCSXc4jwwUUm0zPcNYbCbWsl/LIQe5NmCtaswqjIBc05QRQQE2BaQc0gw
D2hnSFor4TLWOZIKc4+uFmj8DGoMFgWbIS9AiONiNlbEP3rzD32sUt807Fnz+RIo
P2RNU6TFWGVAgplwsWIYU5ullnWs82SHPwhmTESZzySsT5kloMTK9EdfnhNa+r9n
HF8s4SiOlD3UmUIRD0yEeCvHtkDE6NCuzJHNuUx3DrqjiL6iNGRXMphHJgLoZBfE
A2H24XyIlBIWeayT8bEJ60N7Pcers999Hlp31i8jAdMW056MRfulh2AqXCV0lWB1
eskZWxjCnn3GT1Ffe22WiYbjg40a9VaytnQfAMQ7I9JleyRmhX0oiv3Xmah3HKvu
6fnKik16ssr89EF8XmW+0xNpqSg3+NcpKh6YC6BHtQzcZOLkT1NGpzpTc6J5EmRk
e/rx3nJ6Mzuu5nGFVpsy0aQ8orbErGLnWt5Mic7PLSc13Aq+TjPbMAebyyLzmLN+
M4V1UZICqomuXf3UC2o17uMb3QL+5eaTk4BYrbvhiZdi/u0xa1A4q4RHOE2AU0+V
+XwZ9R8+lWVR31R3qLtjoAGKW09suFAK0pW3979gcnHGr7yLOEPzHnyagVHes1iF
KaCzXSu6KSJcPqUSiVlghYB6YLF3q8ofdwBF7P5Z1IzFVzQI7DUfoU2HNjdsGNiF
QlcaA7rKkmDRYI+V4iiJLE5foJVHGHJ4b7kYjedDKwlXTtJ7n8fM3wT0d2zX2kQh
/f7sMuuaxHZ3Jfi1DVibk5NV9nsk2YyhXAYcYg29EUdDQ2E8SoCPPAaVqA9LrH8/
SeTb8qB4gBgFzw+PVl0oH+7SqvEBkbCU3bffqREeBRGtD70cUAnLj/wh32pJtr5o
qs9Gdpj0fg4ud7jW9RwBxjSeOsW32CazZEkNx+24an5a2QfdIGCWQMVO+djsPpUH
1HxGMpHuOz1hcVwHV3OyyXbPZFqRwR1DqoP93GAspd+SNMgyKTPvG919RVEyz3qE
sB5Px0BUOFp5lnCW1nczouUThelQ5iMYMYASAAl5e7ggk77C36f0hGRvpcomydcS
sej/hfLAhGIJurYhhNvrw2h5X39OVdXIftXakvPV0s1jf7+dnElgHpfsUI3QnbQ/
UQjqX4NImN4h7iKSTkL0ynhGW3KwnKDbuKDGQ72AcSv8/xc2iPAPTy6O7qkpR9WZ
yMYcTTXpKUjke79K07xzzVNPF4qP1o6BWPnYywFlOI/OfotkRgcimB9kC6cXbWGa
7Mr7NOmpprRA+Vf4Q3BwDoIpt33tug75GNYRix5pTHmyjVbssLjOMPWCaMFep2Ap
AjuxDrgAq3HxtCH4cWrH2DhdF22JkPFBnDQTe28yx7JZtnGDr0I8oIwuZ+QkoBd/
kY4Rart5O6oPameJ2/7UeiNAfTWZaC93JWyyQWOdTUNaZgznQu5VeFSemXlZSf5u
izNPyO3M719doZa+9R3COWQoVFEizzqOYpReMmH2JFu6lsOyD4Jo3XaTooYcx2oN
9SGoYLz5SXY7tizj5p9hmbmEjO7Zj58JhRm90ypzqHg5zdUYcWqpVg9RGWfFKdV5
C8EH2IRLiBNwdyqeW7FGZq7zQFoGczOpCbOjnq2Yn8SWIqOyWqO0rUodP17rkr4i
D9LoqavZ+yeWwdqaXzBd+3vjx7k8doWEo6pARAW9iTjm1ypjtX1IurqT1hpiAI3d
o2+nbBgaBLQptGPlUShgHp6w1dhFZOLvhsM+aTXFl4T6Uz8U9Q51CS5TGR2KuDkr
jL6EfkacPFIVDDdG9we2TU699NouD7U1REUww9265BSFl7rCUr06nBilIo9QbPdk
laD3zjsp10ZoeVMBVvdwfE9WVaq0xWAYi0MY5zV928J4/UI28eyQf+5Il9H2798x
rARjlejM7HTTQddfjtvqZOtslvN9vAtqxWHt57qDInAN4WohtgHGI7p5YOAPRzl6
zwllOp8/dG9JlAS+5zY/6IvJLpXfZSPJgAA/CkzmEOoEO4gjudEpTk7AZRM85bxj
jaYqxIBSvsHjTO4Q+KfuNqgQ+ziOZisp2ubvra0UHnosw8X97UbunOZjgd2D5rtZ
//pky69hR0a8H0fMKvHiGfOnL/7n30PxwfCRBSAtnfyNQZMTsmemYs3LVDQgThBu
IlWPRKD8ZYqMCAXVRRieLKhcZupF3VHNMSFCUpb3lIrdIz2oCT/hxJc2pQBmRSuM
ZnFHkbbNB2V/DyWvar2IW/pEJbNTTjQuHQoKOuy4+hNF8Ddq52PWPofA3s+0Hjvh
Zu0eS78wiZ8c+xGYt8H3RJr7ryriJ/F06Ynhh4CZ10IMqm0+l02iFHG6UHCJ2Z0Z
9xiaP0VcTHOE0uBiScsOJgZMe2buxWvT0X1J5eckNGVEc5NKeUHr7vODHm9HKZJE
Su8ZXkTdWTIaYgFDrCYx2YjLlsx846q2jm6MUcvwU1IlyiUUYiMB4CwIKc1kj85h
fiJKuwa75IICHKfId1glZh9WhXvTmxXl0E3hEBSGmQWmUY3pmHe92Drbh4PGS94D
bp7kCAFg/21oeNHvB3xKV/yyR2Y5lE9EJLCUTdWuaARPh8P3WWZZVoWgLYBpWG9g
ZPzCZJo70E09F9Qa9k6BIa24vQEoN+kzVuS4r8M+QPSwJ/hT1V+vlWT4QLcPRLiq
OqA6P/1bP1rCYgsHbrqgMmZvCUQj5ofIfJNjAe0jW9rM3KH4FGCHmdJtu9QRHCey
JDY4Q7z/ES0603Bq7GMe/sqytswDZXUEU07SWG+7B4txUMj6cj3PU3YsqFll2ceC
RJbaAFITjSGrAN1T3OfR0TWUymZfBoEeMUe8oeuKf7eWsiWNfGZJx1RiXg3h9KaF
7jU6SCuCuIB93aNtQsdW06LbUoKWX2SDW38+GHbAPuw0cRJB/ZNi5z6wGDP+3zdq
9MOPJNnlRKUZNtusj3sa5eYu984KsrxHBqOW/xxfqjHdbQkdI47nL/dbkeIHH4eS
x+omuUKz12cgO3AkZeyOjALqmBo8WstfmVumC9YufwKU+pGlM8z1dMbF9G/VeVjd
GpFx68Rb+mnE1mrVRNOIUWC2n2IKtCGID7J0tAblpWWJ+30B1FhWZ/VmkrIVDqNC
sWIQxnthgmeMsupnxNMvRsW665/fxc1hle8xTkm1/bGfzzTm9QS2rvJHUJqN7nNG
vzC4sPk/7m4uBMFZFTlMk+UyTyONa93j3dwVNIxIkUGPc4v1SxBs3TX4sdPcCPZD
wgL6ZBg7i/OsIsE0MWGmntU7kZzqDYrSzg9eztV9DSF5fZvmucewAUstLQrY+4Qx
KqFT9FAGX97XEJmaFfD9lOtXPCocUU/PYKh+hmCPMZdst5NGf1gROK0NHKUngHeZ
7he01xR4pN8Ca4izq7aQ68tKokHPPdZ99+ibe+i8fQ08gfrHia912zxqgGXGtt0c
PsFSCsRSSVzYnMCcg7h+vS83QXpb46OPnErO19uNtMGqsGXogtpe/t5bvKt8M7xY
s2hBaIlKEnQoWwzkA5Gx4mkozZTU9MPGQDHyYJibTafbPWoVvGSOv7nRokba6f7i
nuCkKC/M1rrdbh4nMG2BWIv+bPt1kkostXsX1WiN5Wbvb0cksLwZ4vgJGNOz1C0z
I1jHqliBsrdY3E4rYh0Tl949NVXKRSAbZ7dn5cRdrZy0sTbCWnzw8OlbMgK0jY9A
lOz1MayVDoAh2x+0AxWbRBFimGRzV/FoeFa/2dqbgKgmtzWpH2JWf0PsJghnOoqv
cVolfWyQey6GEyQbLzXl0O8scHDjFuXOEF8wivwtVbRxA/TzkdKjjhk20wSD87Zq
mE0y2H6D3PLR1BQo8A6/7VlsncbGR/pXacYp+hklxLYlRBs4aOO21yj3WuGM849P
fvg8AFdGcyC2IxUkFsJoXoJeVzCBRiveMC3dWKg9ttR7MaDPZMUZ1x5J7jlq6RZo
EtWFjEV1FpoOGaeQknA5W/6pBXBnOjtXhYsPWPf9Mm0WyGsJlbHXrfj2kL6dLolN
CgxjMq3vZKmUOaOwsOTlwzD3VWDl/3Gmi0V+tPA5VVp96FVd+7X7LOAjiM63cxa+
tVICnOfN2F1jgitTLuDorrUMLlRsUE4AUHKPzkIbDDEFMbTUm3O1WkVf0TxmN+s0
JjF3y3MZpG8EdSpZpn9T1M5cAyz9h7fk1ts750HBQPUGD22eB72BFkWySj0ZtB+2
i+wByBbcSZkIg/Q2LiOfde8wVIOe0pIh6Q8l49i5syUoc3opd1Cl6sgauLX3divi
2RkGUXdRvJSXYxXdQ7SCdkhNz9A5O8LfQJDjtMy0KHBmJ6BKBaL/HixITwv3SsFz
hUxa2tg0yKbSmc3O38RIF0S97iYH2blKThzpru8JBJWseyYg0NwtvBxupsx8rJTL
EZq0xz2IVgygikXTKPzh2Zq4/ZbklsWLMTs3C6lASGlHIFtZDxAKIQhhVnU+PNFW
0U6fp/PFPxkhPghbt7+bagMqo/+cuDLsiMQFCjvNHhslZZknFdOG27chZ3YHsquX
TWx9yUznXqN96LEDV0r0hEQEuPn8WejCpPdEIO80wUiT+rbNlRLBgVg4NrvTvmnc
k7ET6pETOFWnCroXx7GWducYd5g9DFW5/Xl133KfFIIi/MLZP4RFbS5+pBTo+ZSi
Mfi9uchUm1+fOmovYQMZNyScJyowuwdo+kdO7W+jn1QCdMIDhW7GNdR24uKrbNfy
VRGx9vei8ORYMGkugxh/KgkYnsqQ6wKTHfi76EkgOUif1mX89Wwv9c27iZd02YP1
LZu3j26ue14gInZytU6zWNu4h6FfXa52VUVr/IcppNFuKRtAPXvrDCxFN4tjn+cb
iG1eB42hC1Z2G8dKQUE+DZxY2c2xVBcR54knhsexV+QywxJHeKMc2elv+V2yc4Vl
D4vU9zxgYLZ+dUQ4VvUguiWeDrc5HUEAYAM2ci6jkFASlK6o5Q0/RETqZ10rxeF2
2jvFvr3VZhQGHIb2Fk1uFmt7Jn5Rg46ntYCq57Skhl+d+wIRqewBK6lBU+kZU4oj
LAjc4dxUu65Bw6S/L8mswJ8WYfAM89jFXrMFI6tvCXf3qbCUfAY7gGaK+ntNFaVo
0a3dFNONSeA2lXAX3MXbcF9Ojg4QIy1brZ4FzdnJ+iPzyI92apu2jK1b6hB7uu+f
TH4qT4RFiAuYRDxOh88yvZtq8N+XhBNa1TFbS6m6r55vztj7Ea7i29bDW2Wd/1EQ
gEKvPiiezyBV7z54HtpzjR32SW3cyhm9UoBp3x/TqDoc+RFidHfvoN8n+h3uJWvU
wcDbCdj9TMLyE3R33u0sWyaxPQnfb1JU1+Awik1V6FbNH1YuTO1zCp6xUBHBT73i
lCIBHpsRUhXJ2o/nReLUqzTeSP+Y6S2OAJRdW2RKif/GnsW5dNjAG5uEZrpdkEpF
zVed8qqzRTipxHd8g0VS578f8ByTVO4E2EWWRB0RkOKcwcum60PlqUQFA61uz9bd
BAOd4OvXdqehPr00pLeNuzv0oAqlJchPOI9Wn+dgm1skGOQT3WoRXbb5EFCYYuKx
oSs/nLy1YgdOLzGyI05ftkSA2EWPi4f65KjGnYOtNeOq9eXkjTYjK4fQXaoMoxZi
sznhLUo8GFsEwkbEbTmNvTHsq0h/zcJS4fJs6j31AozNKlCEvJ5jPaZfg7ivcioJ
gTe+kwAL9kHQSKOsTWicZCPAmHxGFKitxrHaXL3nSViZbLVJq6zCwXWj1ryxWM3L
nbptc5ebvTifbVAYXDQIC7p59VOiIvbLWpE5pDFWkK+0MyUQv/cWWtupzG72s0u2
Fce29lFdzwZd7rQ5/K32+p8QNWuP8eF9Jrw0dKSZv7+4BsHCJO0CDrvHNwVTeAy7
YCii6qSVTDnSnflFj3KrAZTJZQ1O/WDBMAE0odRvDRsO+E8BmGw2N6sgIFrbZmCC
wr2EI89UVUIBvEsNX3ME85BahrSIvqosqlZmszFmeb8zkwlVHizRA/J/1a6sA1Wg
r4Y59H+wxkyGE4AwVY/+8rvfACtzA1Xd1HHZ56Ij/XMFlgf6qBcIZu3cpBNf6Qcb
Lk+qaEuT0xlerJrRc3mSwt3/ChQJ+dvLhZCfr8s1LdYLvWGtkEedRKb6PTmQNSSy
1+SFw/GzxX1+GBLphFRtYmRltuHJMGqt7cfzs7+9Mzc7ABSDQYCqvUv4FuMD4LJD
lQGhb6aa5pNBZTAf5b2pHF5GbJivL+ruzJgWMkhb+KAMlbfG7JT1rDX4Acxyt+qW
EkYQn2jXlUJh7z2M50fla/M7tlAl8MifshZQc/Jzd9oa4TnMjuv87RhxPsFethhl
nZTk39Pt9GN6lQcdwsunYkwnXzXipl7QF/NtvWPQJOjy1hdRtMNDjvEdH5O/GVVK
5Hm0S/46wAWy5z3b6bhpDxYFLMJG1QJqPmU1P+G4OjxqQ8+TBC5tVEwKy8tuAB2q
u9eyhjM/XudHUaayZKdvyuAopKznT8p83vd79gJGdgFMWTkI/KhGcBt934ddKJRW
4vf9itnEOgcXFN6dvl6wqElACH22FDGfuaDRRWopk3TSDuFRkxBY32rZMkGCeBF9
BPcxPCBB3RUvYabDRgNapz2n/EW3TV73+6YC7HJXAEfrw3wQN/28gLs24mfrQLsx
TwiRqQBK/vFjugejQYFYvZikrVOjDndsz9Xi2eHXjUsrGfjnQrKQtE3G6AnDvKar
GqLYzegwrqWgLp+HMipLllfxC1loBt8agb1zIUYN8/G/AIe+h5kXVHpLTjCC/zFU
zFYoS7GNkn7w21F2Yaro0IZRWIxEGV9qIPJmiCeixRseeD8cSWa0+hVOMQVh9jkT
p7b3WK/IrG6FgIwMOAKruWAIGk+32KqXzCUV2l1c5PgcWuNp+sSq/LkXfIwnfUF0
agQR0R12HckEeeNFRCO3Bx4XkqqK0l7NUqoRnFhRjTVkc7eAeH6J//rZUfjebjQZ
LqkY/o3t1oWYxswkRir3aBjGNBze8LwCHq+5xEdCmwso2YdviQTGJctutbj9sTss
Mmr7yvxlt8qaAPFQjLvGwcMxc/k2A6ONTqj8rgWJ9HqmV+PUqN+AzS8VabUPleQw
tkdJEZpfqL0FJsZ9WtwItetj5mx51me6ikC6YLHUcXJDagRFt9oowZdVxzd65A77
CD0B49Z50T51Cp/Q9cDTVm2/JyNDgzazq4SDM99NPoFkmIUl9/pFK4QKRDJ/XJdO
gQ6C14JRQDvLxQO13S4gF3ZwFGgyjmmeZdZL+UHhpJJK/4qIdu0UWsbCC+IO/oM2
CRr60A0h+eta5nRuJXNeBeidzg51Umhj9T0301hYppb5ncYdwYRBGfb3NUqjaOzD
SFa8FSSs5VxvwkLx+W7vpOt3DMfmm0wOzR5cnm2l0i0E/sEsaaGAe4QpE9iGjpcg
JYaPRONvQVh/D0cWoghOyjgsJMgrNkxDmwdynyNKla2mleb0+hAUye8cFyFfe06N
wGBW76I+TZc0AGnDHniY/BCH9x8xyIDY2XJhIugYZckS3iOKnoZ/uTcci4PigBy0
1SLjZnBKhxEJIAhgmZX9zWEfWsd3cry7+e65ll4iuWSI4fTqOTdZGu+AJppWcL7w
eqdna7SJHnLVeeCo6FRv0/A2grigXigvcIxgYBmU+gfrqvrv6GgPrGejPl0IvMPl
WdwvZhK1dljm9M+8tQsCs/yu9bQQ9iuRn45x5FWH5x6EzL3nA3XacDbvYB3QG/3+
uM2/6fsZTB23IsaDl9Wz+n1jNXBQPMfHOj9di1iPO7Pu6v1WJdn67CTRFUyjMvWw
DOAWzNXxdo1ltHl1EZXEhvTwOd5OB19za5IfPfaw/wdZZKqp6I8JkqzlwLcB2CwV
WiT5N/+lEMhr8OFahlzbQOX1kZnMwxIQzY4j61lbjDUFpxZD9/Rye6qVaL1RgCv2
NRaeOtuOLZ0gUxsuHgeWhQuBZRhd/P5hWhaO6tuNy0zNLtkwzn5ydu8ORlBiS7At
pLiA2yoDTLfl2q52WN994GNROUElfc58n2C/h+mLFExfaH05CxZynp5ntAWfz/Xw
QzwjWob0VvcKa9fjDXsIbcLUBiMZNoPTVjxV6JDTbq6hoJwMq3IA6yiLntfZBIU8
wAsrHSHovbPiugZufbAnU5uWoszRL9PcfWt5Lf/MEyNiaMmtJwQ244Mzf74F/lH1
XibRrgKI4qWS88I/vNt0NHOCDNf+DLkdHHp7X/0++xRQlvbaLkHTFoy3D3fRqgBU
vGkt6qyQKlSYs5UE12mxOvjQnnHMxN50HK3ZmQnj2uwqgZA6qCzLNcpAykuir1bU
fCks6V+9WXzSOEFkPNrQs+IuVKdiZYogodnT9rsKZ4X+McGVoikHt3Ay9oJ3aVNI
cuymj5GziZ9BczJMMuWtukeBRN5Gqm2LbOgOajtfn1CrPOG1NpDtDPNgTHvXv852
GFOFvq9MmnHJLk8FXp00r46NBmQKDj2rPQWoeBJSh5oD2WTwsyMxFNtey8PiBu9h
3lU4UrSrX7EEGa+aFFBfri3KKJU0+KeEOGU4BhZ/S51A1nbvQUhHpOUjk0LwuhLf
AM+9ApRcNed4XPJJKjCRKFu10WA0O2C3SZhPquEwpn8YdT9gkszHVK3IiakIA51l
3KBsv8FsV+tcX3f507SJNx2e0l8YaY0oLu1Zp1lHEvF4CckEYb47e6MT0jHaDXU5
umDlLyDPeQYIx9apLuhKNjNlsz0IE7ZcMMMXWkmZwZJ0FRmpCsKRojx2eVF8RUmb
Wu52Kr6L4v/qm43kQiqTrNLrhvulsrRliCSyFATBkwX17ULsSxWmbi2ttBhx8xBz
NqEPMjz5gJplXzOdPF5OM/ughn0WwXM9ixl8gU37Pegs0wTx9RcepH30ZmDbzlPn
g6DLfNVQ/5wF0vsW0g+kx/i+quKcnoDDjCB3I98D42LWAk1Kt5k2qysKIzIAJF2s
0779LIuQNqYsP7aoDbqXnW9NKUGeGnhNSaglCgZZiUKEWzVtHrVxTLeZCwvZVptK
jU3JlOdgp/Kn47T8TJVIr88pFwCOKAWD8pBWR9ovtKl0RJ7TaRROVAXP7krQMvYs
TEH93h8tdWFRyTCCmKRqUPosMV0O6vJIv8W76Jx1xyuCIxG5WcN+1z4L1dkYDgl0
kOEJngPNDsJs/0o+X9JoYwtDN2BR7WsZ0jOVTkGwV1BIQ/T2E3s8uJsdZK/ddSqU
fUg6Ge8dBIxYEw7YqpgCU06tYcgeP4bGwMa0wt0ltNRME5xihYdccS8/rzaoKlpF
5pQeg5qft1orx3ipCgtllwhn4iWHRjw5Mo/xJw6+kaDE8R/BrjjnrKZG8nKZtzNI
S2QkhjL/INOCkE2VHmOxxJI3sKUXkYQvSxOJbS5rbXPJm4iRRiMHZQoKn3imkMGI
kxuGOXDBFPNI6B2SNL7owWl+89OTgjde8HEez6Tam/hUooziLBDo5Gkp33FICNU9
kTjvLvLEq55UikP0VNWNur7rsbWsMW7gMvTprgVq1wYspQ+N1zQFTHQeXyw7PkuG
UdBuRinIn3iL0rBHxltYdOxza4U7/ZPqyh76/Y+JBEKN2qX+/gFhbgDyTcvFom2M
oLn3nMTYUKtq2KYEKBDUPL14OM/EPdaAHX9gDfZvyK+CQYjhBM2xdIOXyPNdcqwv
1aQ+Yu6PB+GgeXHm5phqbn98HW/qlYFqviREfm7nFJ47HcQNcbUVpJWWPLGIm12k
tCeEr/BBw12GNmBpoB1P8wVv9hmzasYfF5pkctDajBzjUz9WiNxASL2N9hb/wDW/
o3VGL0TxdSKijAIsozi753CzqRxecTWJ5gqytj5gsNBpOUFx7Uk7hNbKIbSg153B
ywA9M9PtG3fWBDSNHrtbfsCGzVwMFkQdaB0+i/CdqTZyQZRUiIsw2wRAlbF2aE8q
Tl1aHyQad/0LQRHpb9uuMoWnSrIsy/PxMOBItVfjKJNrR673uBMo58RKl5Yucp4U
rMCRgA4cf3pFOgYVs92WcV6gue7CQhkzOMYbtElQFz36h2DOsQKQaJ2PkTxTUvP4
WIdpRY//Aj7/j9+q4niewlffLfgoW7N1PEptUC5CYnJYKJpmixTfNoKdAtsrwQno
qvjsDN9mFpbukgh+wLoQg4OAUdpz5DLb81g54DtW2scEm1tQrwguu4RdeUB3xISI
OuBJtohpDAD5zVGTpWWUBCnWNI62BaVG6PMJ84ng7oYPYN7rhnM1VsFBnAX1C/PK
K6OM+Nq2YNGbDJJeKkqaurLbEH+ikeekxAbr2UhBJGzWEHLosYGzGVwG51QRWobW
oaTW2pRhE0QobGCuKR2DqwOjmLSr7hwRIREYDH3KyK1h7mQhk3+gi2lgdBZZMhTW
DeJ9O46ELTKSvkdNMaDtQWHDIYmx8Nz9asqvSJEY0l4cNUZek8JJ7ukNWTMwLtha
h4vx+ii6qwN3x9TyIitcROjvXiOuMYM5JNWWoTze6s1PwtcrFtmdpU0MybBGmZg8
/yK2HPdD+QaFz9mb4zWOTL2drB/DyGt8JnTuwsa4HAwCeVgkgnkYTaRBjQ5OX0Yc
bJKUZY0rRsjb1oMBXGNLaZQOWlTdZ6kBQtabA5//T9Z17cqVT4gcpCpwicRENkmG
JLeaEBddSbR6amdO5x0a/wUnwl48AWOojzroRetaTOw0wgsSR+tfuwRufOmQKYvk
kt5CIGuYnxdE2s3sraeRUvmPQmZA436HmKnxeMOlZwVsp8T5+gK9dzevkYBeRVX0
pNU4lbWOMQgYziighKtZsLXBZzofzTW9WArG4sSl94sYFftMBbWh7m2q/JhuspHV
KMw4J98VhURPGIElJoYisNE0KaPP0nnYKCc1hKibIYCvkuBi51Our7GcG7KPTjU6
RoNWimRdyI9L3dOL0lU7MboIjAdXsVS3395VUfmysBP/fSzkUJj0chMtVEUnTBad
KxeLz93Dy4xzsmNTtsX1aaNqbNE7cLEAyxPPfxE1xKUKNK5vGVUWi+jcwUDeDOm7
TI9/DpXBmL1wSopJqIojoPR0HKG+M5E34ha+qgebjF3DEBtdK0NnJ/gfwthB1gxH
OIt7cxxY+f8Q2wO2M/7rU0zyaDsS+f8ZWdLZ+6Vh9bBZ0G2dddhtUWnpumb7Np6w
D3OBrg2on29yoom0GxcbgIM561/oMJakd1Q/ZtT9CNwIfDl8bNjkGvHPM8l/iYzM
GbbQHzfKHlZJu3jp9KL/2Gv3s4v+3iLxb++6BkSZ73+bCZdQ0Eo6aaLkwWjXvU9T
H9c40G4KioNan01jfspseH3MVIaWl43SjQoMHAXxyDO6wJXuckeo2yb66am9Wy10
A1EUrBb5aajNbKr2KforWLt3wF98vrVPG6aV5w9ByFDXx2dv86YYZvvirOr6Vs5q
EWSmy1tBQAMk0ZWknX0dfpVLfJEmGSNotckEYbmGD0Alh9kPlhV1ukQ7IMt60YNJ
osdf3i5GZruNfPR+86i/799i+NiPBE6E5DWzrmc9lZ5XMUGmxIfsybYW3nvbVvlf
kTQW7dfA/ftk8Rue8btUV8DUTN04pPAu3xYbrq/A8Ak58IEF+DSmaa67k0haTzkI
X9k3cHbNxAwMyDgHekhx5tW5E/Z2lVcgvBd7rywGeSpLFpl6ipy/kxGSHToQ1zZ3
NCljheiunPbgXANJXss0jpt3sJ6W/tYwJKbqWUghcIS9PJWuXE9YZPYm012Sql9E
av6SfTo4II2ZyxoXj45McnB9ldPYjamXVXt+23jIiRnZ9KlsrjXcmx0wsx/ZnzMd
M5KruafxACd0MTFOfOkY8+QhLVj2LY1Yb4fEwOeUW8ATbCGCjVd5gC1CZSW0jxnL
drTG93KsM8g23X3KBzLrBA7epRe120iymckbafPQDyYpkxiEUM7KdRSOhd4y8Wyv
0jrluJVqz9iizmD/vjlAinkDzWe1EPQ8V9wl6+rYtKa/YOve72PHDpICdwWRpn57
Ji+5aiAmFHT1v1YAHkJnV2WoAatr7SJ0eUq9Q+3Eqz8DOJPrLV73E+ljMx2dGVlu
CHmBr6sF2jFNBWP5AfcuGs5dM7Dj8S57q3K2iplfMhWzTQKzDPLAdXXGULDdUyWX
xF6yjO3J1u8uFIqh8Er8ZU1AHL1ZbMD66ydUzO7jHUPF6TZ2dlG8Jh3bdGaAwl0x
HCvl1ch6X6W5lR2dfRLeJ6JyxmdNUSv9+cUKn2GN5Et+iOnvtG/4pg1l0nA4CVE7
0BplbVuIJbQPuYtggvfG5yKzTHO48x9VAMQPaTRb69wRZ312TPypTMK+BWVnoAJX
2Q1LOiNcxthS4waXcF30T0eEsBTIj1jIO3z74g1i363tbKrjtb8QbeSch4Y0lhpZ
JL3IQZTPoSnygnlu2dAZZrX4Kb2OTJOAqJMvIJk0AKzlU+4d0hsNTEg0E9qKJtXV
eroY+ByREg4tIDvku/S7f/w4WiQF5e0l2a2lNceipmXu5WYyYo4jC5VTuGnvjnS9
mTpas46Z7Q4pzI8ipYzRkWgm4yplbw2x90rVxI3tAyxQsCeSFRH2Na/hWtKc8Nyx
zZZJmd6+NzXvCnPmnU5eCNejTroE+YXvDsV2/feG5Bw9+ePSSbfc5Aaoi7n9oGvF
rHF0F8J4mRedSXp1yqdi7TcfIcmKKRHgEQYqJbJQZzDrXYZzqIxNrf8CrG6rRH59
7G35KkRCcGD6JY/CTL4upg18ZJjW3EAbAsyoJPof4Dn+3XFGc8tkmtAFcmFILUuv
elZ1r9ho+MvNx0W+ePyaSxxYD5ElUYrgKjcQzkcLhpVN2jEVsl4E0Z5vzeNMBoXK
VKrLndwnvVDaAg1ePY5cjgFoLIzkf6fCT8fx+9zZBtw18IkH1H6Zm7jEUAlw0m5x
NskySwDebfDCfguCTQcBSdwnmVuSE8LLhQJLJyV7M9gdmVm2gc/Xzf8IDju1tYUk
rXT+fpSrAf7eB7ZjeQ3J8GW3xrQrLPIPGY2Tj2gcW2nD213jgjbPxx1EXY/2IMkh
ar+pIUwRnEQRyUPFtPD4JWxTYl35xVQv1o5u0v8YpiDTm3ZiG6swTKCH/5noeMv5
Biprsg30f/FXm/I5C9LmW2Rl0ItEWoptiwksl8uv8iEtFWbw9JEk29dybPO1c7Nu
aDLyTTAMF6BfZAaVpDz8dlWMRLyPWAvPKP2eGCesbx7vMuDyiK63y/aRUtP2PS/c
nCyxEQpeExSpzOkJskgnHwYhtj76FcIUlkQ/ZoLcCO/j/jGDobncNeF9aRvQrL+P
te/dzGc8EAwRYsZ0NDc0CQJZ3UfxcRYdamvTXYqRvVUbgdHFeImHvMpuwRtgVrbz
MkDMQPHOhHKbRCMuthwTZoF3gX4q9gL6t/swKb7gGd6o6w7MVxfX+g6xufLSe4V/
9dRtvcWolqqL8OXrwoa5Lsk1a6tZgSmnXws5SX9vtkwjFYwUXnRruQhnmN0vsDKy
KAE9kDCB+/PsFTp++HoaSNoedeOnm0qTO5+6mfpBr314uX659xZMzcs8Q5bDVM6r
xIWpE8g99Vr1Z52MuPkDpi86Gwla9OUupgST9a0ruRyDaMQ12/ka9CdGLJTQ9hU+
cutF2WEOrWW85qqoOpTmhhD+YGhDpVW5E1xWZStDT1WlHeI7gLc6ICmTGGOmkrdY
xxQUPv63woYx5DBi7JbCRkbnwLn5X/PRWl3bUAAP6ssfNfl2CLOslu4iPtKzW22y
q8GkghhujWh48MdbtqVi3UjCrpK4sI/48OvDI6PNlnunXNPaBVuFm1IhPCDpdc3s
IPtVcXWk2b3KbPSOK7BDvjyskcdlb70u8bOTigs8IFVsVdZ9pmF8Y4KHLQuXXVe9
+0dJmCGCkGA5uEKQml2h0HJojuIH5q+e4UOjC+fx3gaE9f0oOR2Kd7Y8bGnqvg7c
BbldCmrHuIN2K45n3n11TlrKTTsdYD832eEwEZTwFz/gdur1TPbXltsrMvN9/ggM
QHQm6ARHfXgpt5T2FJPbj85ry/FiqQNSj7VAhVn55qj3o70jAbYPxX/iHGee/iY+
rOYiQ52FV3lN0H2RFavuK+/1EpFciehwpoejYIOny7wfnesbylf6ycVDaZvjTm1y
ilru5ggrzb3TQAAbF/b1Nb61r/ex5aUnivBPbWtySxmyiViIAYU5wVBb44E00JVq
LkXJvKV7SklBe1BIEvteJ7+KbLLZjlJOlnUZRQwAlqMSowWjKt/2fZ/Kr/ApgC4/
MmL3iwdDuGUjotLZ08TMt9YnQHxw8aV9l6bB6cSl3WEXg92AviwnjK6vFy5Ik7sS
HUvq6DjAIiA6kWwKY2eHdrCfEiw0bbHhmk3NO/8hWDKNpYheBS1JGMjEBP+QsGGA
lKMLdj0hXGNBaTvap6Dggmz5VMUJqnjdtStH4FUefKU1zZs0WATA4OifgyJokSV1
TGsURWGAB2Libgc+HFg4WHBhQ1aZPDwpvhh6WO8yDHX+eTgKg9gd1EEBqQkoWsc0
cx7VLSQ1AUawhC9zuldgbUHe+vIG1g25wXfGzXbZzs1zisw5ZX6O1qMpveGEaVgO
dU6UPnUCX1oBOFcw+Y2Dtz3zUakq0tDYELRS/wSiNjDfWy6Rno1DrwTDUMYSR5NA
MtwNzlK5S7JW6bs6nu3ooiV2YrwCNAsnC16tNyzwF+inig3sMmgEA2ODs8h8h8v5
jQz5ztaR8oHcdBIJIVAilSrW2umOI0+FT34Na6LspMc6YwGms7edAmu3U0QqcaaO
egZAN4AlfctTxhC/EYCRYfg15SRBWDtIetPo6mOEIIRRt28gBuf8m3Xf2NdWMPzp
D5pBQqoJBphy0/TanvXPuEy3E7ev+H3KtaCbgAcrSTR/ZkzUSMZ/9OQhq6s20sWW
hohRMToJe8tMgve6Oybm8TANSX8uiu7VQbElxfuPlRxfhhumUPVahnPQdj5sCC6a
E+u/IwbvxX9SiUF4/0avTGmD3l4SYUeAIcaR8Hm+1TVKOoKVXx5HFS033ju/i43X
kEJo3dtxfkKXy3U38dgh3iBXl7saxe+yZJriA8xGvARbkc9zqaIOoE4s4nl7cxVV
hV0HbPtBh5pjYJowC6IT7KUR6EMgj2vpVId9FXJhaxbsOdBeBT8DWmKfwo27T6W/
5qNfp6YYwVdhKrsBRnMZJZRCeFQa8NPEOIkmRM2Mg6maZMLshPvF/waa5xK7KUog
VAbZ5jV51Uh8RMu2aoAJrSz7jvi+ch4fCublO0UCa2rLq3HtJSw/Q4pRarp0LGTE
Y6tnRyizRLAow0YOMS024Qr/ORIaG1DngoY4go+Nf1CehkQ3Ob1yc+v7P8DiMqQi
W51KsR7Y5p1a9viMcb2/QAU05uwLwipht+Fwoc3BOTIE2hnPC6ZOIhsVV3FyPYDO
31p+VO99DaY8WZqg5S6CtJO8uIQGOIy9xIL/+GjlSs+5L1TI5HuMH5YysHoZtU6R
YMlxQE38W92kNvZiL3Gtsp1MWCYNazgtQBITBL0m6OKUIUaCMeu7qpzFh6HO9HC1
Hlm6rxOhBLf/+OPauJCmybdxaPDAakRURFGiCGnhhA3iF8pmkp/f/Pxlm+A0dk9e
5wW0yyrz0TbQfnjz87J16wdxQWZ+ld56j7k2oPM6sQ3QEvsoWEGAFqZ8IeQkM4YB
1jg1xtjlhzziEB12G0rm8iP4Ty5wzDSip0XsY2qhmwo2gOwJNCqe87vrm65MOtFw
i0ea+EQ43W1B6Ybw8NGXd3q/v12jDHu9KbeCanqZr7opXQfi5OahOpJ6LlqDqDgV
qFA2YxogXhxKiZH8687qteONnmcl2JNi2NzRfnBT72BMktUktLEKns+gSAvVjumV
22rmepkwzhrJOPQxVXocHLc46rzQc9uONfYMxrJxSuLiuVQnY4wgVP+AzgElbDGX
vs4Qc5wLrndl6ihK49PqQR+ijWw6mT8Cxi6MzvcVh6hRvFYzMElS0d7HrNfgbfhs
lMD+h5F9MukT+3a4OAuT0FX6mRIZJp0DbEjIi9c32XZoC5g4Zc1KEi+DpwWFh8W2
kNR/f8iwvnZ6d/mWlCYWz+bYZVogyzUX9l59MPnb7oaV7MIn3lIeogMJoldVDuJf
oRFOQiy1Z7mjHy+RvI64ZlcQBvyTbJdXrnX/J9FdNNYxHmWHbmQUKa7Jr5v4kNYg
HANbNevo1YjHdNE4d3nVpemv4o7Yuj4DXpi0dJbV4z7FL6ZPE7TpSyLHGEjUlxh6
sqaTM1AbNm9u4PJRnu4sJXvY3cQhhD3NsLT0wGulBPIYZmlRJY0Uvf13SdUhRI2F
vN+P0mTgrZkNpe65YGrXZIcS8Bx93nN+V78bHq2SW+NmPdG02EuNIqAvcJhCj6jc
+5iWHOwOCuCnjnUBD1B1MzHx7TTC3w23MF7aRotjI2ytuNEKqThkseX40NK4nC4R
xR5ht1J1pNL399OesvcgNDTKuN7wF3ZgdKTvdge3DIdMtWMVgKIu1AugbH1ooQx0
/uAHI1wqn6A4JeJQ3X+/2UHO8SHXeR/kus5o/YpN7AD/5q/hjQdhBIT2K+7DKxL1
yfLQvPgbjaPV1mO5zmlkyPE1TX4fY+KszoJKxcppfU/D68mhCchlxbBrIiXwgvuO
sJMa6cqtBvRxEA/BMn5eerk4cufLMWdI5McMHRgWKqgd/5q6seTsJxVNHVwnOoHq
4OPxuR5XZg7TO2ZWS1JoYBsyQY4RBSb+KsAr2pIqLSbzykDCEI3UmcY58d8nuSOF
ZLpApEMAARVXzgI+8Yb2OMDnoInmbsJJosmDq56h9JmD9pM/SUvinhyZr64rMhUF
UyZ0AxgSqFYK+4gGzkMG2i6rIkQCOEhLhAkHCJCrVoHCsqqRfxyO7kOrRui0oCO6
PJOzw8Pkl5I9WqrToAprzrY1FMyTUqNa43uOCZeHm97D8uHTlb9B9U8bxy0q6ZHL
LnFDLlD/QtwENJYoLIHUAYH5QSGHZYuzmZ8+j5FFBvO8dSYFKRsm0FDsNI15oeqQ
95sk84ntux6gTqseztxu4Nh037XpSpDlEY/nxbYFx4YDLSGJ4OoPBIH2IpC86Fu0
/pdqJ1uWsDTFNOWvVC//iGbsKWdCdaE4CZ+mGt/epKOg9Fa8YG2AyC4/nXtIwPfZ
2F1Lne2Qbtwc87XO+U7NBMzxQlPJso57VirjbbxyWsbBL+0hyooeON+V0tt9twMM
lGUyQ3PhKs183Gxoz9Fl7DDUkFszlZ0whUggyWnhjc8EFBHrGN9bmFsrSmyKgeRH
Hzb6gQ1lOFpsrpdu7PP/6PiLHpVuaODjRkvrSplBiMuUiJ84PULZH9Hz4/cr5jtY
I49vEZk1UXTvFSviQXn0Gvvg64H4bflCuuH3v/4pEn3kNClSoJwcu8fVhQBt3I9e
w86g1XkNTwDzK7iQult+c4wFUcJoTe2I4TGk4f1qe/F7jWPlVgKigBo4nn2WvsWf
+mhMmqAk+rE91uAysOph+5NrEyf/ZxH0Xc18AUl23WqfdjtAZO2btEQUj18q2jwd
hAtGCbcjZN99XOIG5lkZwnXrw5c5kNxOmhU8svfvC5jssyMKtutfM1/8t1auHv0b
PHWtHKByMOXsp7X3JRn3HA6NIjF10JDZnff/MhgMStFIY/CPeLgf5LBQ+rHQUKqc
g0NZIagtO4YzA0MiYxr6xJAnz0wEqkAwcIUeiUpVJTwyYHGndl8Vm/38jbSd2Q7b
TIRva2p+h7WkXypsqCIVg7PW+r/p0X1OIPiJOTKSfKpkMSRoU7RDnRc0xmIlPkJf
8A3efpb3oO4/2KemXvV8U4fX9EOJhcz61rrhLZQm1NoZxKoaikWt27dc1euaCBN6
yavJ5vwslrm25mOZs+Igsy0LZKFsIi0EuOwKXrf+7Fl8leB63S+tmQ2aT9CbwDY2
UvDI5RlxjbxCpp+vJ5yfI2OSwiKz83zX/ByHx0RClndNq5+VwkBTJk+YGLp6cJqF
MxwjbVfNFsPCBqWtOHgR6DYIS1wNM7fcJclDoDIkHmXIquUvGEILb5MyvmVuQihC
y7t1faZxayLTp78QKbEAztL1bKpikLz8CyRsJ3U/p5LDLpK9vQYhRDUGTmnibWuT
rvE/lzvIhd4JVlvE+qO8I0+qyiPV2ET7pjmjcCekT1ZRZ4RGnvCGroHY6BQGeEJM
hkY6onlcyOTOr4s4C+GRvR75gUBmjgBF2E5nkgzA0sB8+VPq7Lc+OMkmI5dvtoPX
zToD2ZF0JaTtuGzYr0jqANA1CfrfvXzfDW+uGU8AFQmmSfNqua0/6bggNKMI6EsV
Mu4JCItpnynVaVyPC+wvZUud8cJ0X5rQdYGGAJyW0D6ZqkkvG2fi4qoaxoubB1mb
H9JhU7F7Crfk7+7oomZqJbNX24Z6s1peX7sqAvwLgKaI+Q51r8vbOO+8AGF0MTkZ
RBBgYmDVl/2tWdW9PLzFCI6nn7VpHODCWFUZLge7UNKad+2ZqdzspVVBoCc+Asno
bk35zd3HXzoxIvOJrJ90uJ+ce+LoItPcCc0GZwdAY9Tnf2geZr8U4eBKAGW6XCPF
GWm2AAjlupqSKWUbBL2myAyM8p6mchbkkduWi1Z5ZaHHN19m4VXwAw6eZ6lD23oJ
FP+J8p15/Vmr95Nc8HuhAr1eY36qLgGx4xozYBEIY0AG2JVmW/qwdDV9YHrf/eRT
i7RK+gi7a+wOex/K1wwNfg/ubChLgUmaJ9+pmYJ0NJ3yBrUNuIqS0xbXmB/ZpQZS
PU9KvHJjLmI1Lq/OZwjRibrVP8D+mQDw8rlsm+4qtM19NCpJbd8iDNMkJ4ouHjyZ
4h2nloMkIKpIxZ1BMy85llvYvD6G/C4adVA0UK3YFHy2QUA7EwV2JgaoStcBX6K7
flx6rLBjyvepbMkP80fMi8blFqtz1qSi9jceelhKQK0jvhRPC8+DeAmWYQugt5yg
n2ScaKvlFsKiWYa5SyF6xu4ed2Qpisxj+kAKoqti6xSZWMhGlWsplPvlx0TV4Sax
lWSFWuSUpfjxr1NcmF39MTZCjOidpDn07hBzRTgpaYlCjoAWy3BzNFtasYLwUUxX
CXkM1sphe7q6dQ89Sffn5KrYjiuQI9rdzk8dbD16TtkWfERuTEz9P+P+S3E0b0vM
EqBRklRjM4CNKBRIK+WzBJud5+gh5yi+MReZD3fnfnu9IgTdxS3qQ7S5cxwTKUWc
5pmvowBKP2x5hr01Pbnbllx8pZqTyVm5/zqwGgnEXmzfF9IE/DCext+4B0DnOXKW
b8r6Euc5XGeoiAf5LhQCSy4onxsE1DUiXEK5+UkSysYsQGa2lJQwlU7OLI3JB3f/
7TeUgwYGE6Z3NyqMAWYajeXgbszUFrq01WPrhg7hIkRmBwqs73zfpbhOB6u2MgUx
bPx9lsORa03CHB5mRN7pvR0lpE1iruuat41/UiL6zuEZKZEmtxVWI2T2LUz7mHIk
txMQ5qTtK+VqAwGC9t65JVEwT0g6m8VynHO0uwhymjHd1scM/DS+MNNOxutmreea
lyzYvgdjxnWjKp6xYB0BWI8X589PV5sW1ia3TPoh+z+wkjs5BGgrYGmBwPTKEZP5
6L8nVDiWrt5gKvxS1Nf/X1bsDu8iOZgZMqnsoq3d/632A2XUEMym1gNBwsSoMp0L
XjwYlr/jbvQsiTXeMyzJdkYfOWffBWlUMzGgaC3B+0RtaqGqR7tcI4i1nbL3cC1s
2CNEdEboQrQbLydBO3D5FWC8mLxc5wVR0KFLcuCiWbmjT2tZcgh4w0UVVTR4EKbP
hjRUQ8BztpfFKVeMSikQgTHpuBx7h5Z5DukqiETdnS0/ly43AHvm/e5cqF6E9+/x
JuJWm8+J1DPSnmoxhTKfgDIGwbmqriTqWldgtS+lJH/CxYIudKvVuneUC8kNz90c
OgzLFmteBYCkQRrcrRJurxsb93qsiz7XwhdMDAjInfhEcBuCSkca+d/XTnCGXk5c
SeobQ4VIEfWYZu+gQD7w9DAX6d1ThovcPN6mN0xuMr0ptiNGcPjquKzleO+6pMgK
4s+fPBxJOYu5RrJvpTfiE8MGLPiAOJQMV+6DTROqZiEgyrrNIfj9yMhbZ8JYjixx
qyHDrWB8HbOqKf3wTkI+dxzfjtQGC3Y35vtrbMlov9tmj2SChxUkuPd5tADIM9Ga
kWWSSnIrUKynfFhsQrHGvVx7qwCXykJrr4ZidgBBHt0zSvgEc0fHBDu9dUHsCD9H
xf+g0qm1adRmaVrExXIjgs8cKqc57ZZdVXyQNlwdDIKb57tsR/c75arUqxT1CUY0
IsqWIjKwwRMW7/O5ga5zKyGiSd+rEj2t7SDD2LMjbM+Nn2KV/jjdbhtx5fC1X+YG
djXTOGRF2plj6wYc5Tx3L1nJLwdTkwFkBwFXzZWNyOrGxK54cEY3jLyP/Y1mXcax
Z4OCuhRvI8Iw9k9GtJz8un47icyNC6EwldZPdpm8elJF/skmUCqJy4luF/zs5Af4
1phbE1xmJxl2h28PFbKYkv9E6O+nZXzYjAJ4lf0yDwmlw1Iy7L7dEIN+X0CMhMI3
Md18eSxraW2Wsdmir3Z+O+FoVjbzUIP308I9yaHi9fhqL55x1FA5Wx49DlI05ao/
YAJ7w8fHKK3Wh7eDN6Jj4ei7Hctdyl9uZpsuOOp/QqcpVd08xseFVXc1L7EXXB3D
xkHhWqQ5qQBXFq48MwkhXWBak115SLvouoDEBPAKtu70GCCxNcjBKfS9AzLhZo1f
i8PWqZFsphWyjH05jHiu3VeXm2rRgaTJfLg+5VJh2ZXSq2lT3AJGj5X7Ek14ejf9
R8R8N6X5WJZ8ZV4qCuXtsKIa6n+S5PH+L2IJ+m0bvOgOEXTUllo+Znrzo5CgcStv
3PCu2GRFylxRbvMF9X4sOYHBadqf8XafMhDpApesK6fx+OBg9voGl3HAeznjx9X8
gi8Y5EVURpC/22yTgoMBwcgPj9RGIWy6WFGR3e9EdPjbxOArnPmjasAD3hKoMb3l
4NjzlL8O3qnAujXFqkS/Ux2GiBqFKo4bL2mMTyFCpUPTE/+u6iR1xXFATx1SH6dS
pXlw6BQakexgt/UzPw6e3qGcj+v7wW9fpSf7QTlAA+RnM1SyFQPVEUGV6fxCHR/d
rGEivZvtVtWWJeUHD7rGkLTJRFnJa3K551Y59A3ccO/4HfziPaUIZieyujxL5WxX
eioFoyPzAUZG7QLT2oJvgHWKeSxiol4+/4lStI4Of5Hh5b2FzmpR4CgyS9AWBKcB
WZ7NHwREse60fvbT8+eINuzQx5wuKmUUZLaUAs00cbGjcUIlvc+61xaMmoucFoaN
v7PHmGVdiBnAGM9ooVCqQ2w+yMh5gMWaPyP6mR0ii5Rad6fGx/wr2PBbHTEQ6DY1
jBuSF5oiX4UVdRBXh/FB0VTChO1FeIHVxlTmJ5ceMVokO+vMZ4954D36RHlMlRmc
NYYIjgRgqall+gISejp3xmfZ/BJzSJhBJ1wYXYvLjrWEoTHxhxszoMo5alUCrOyK
2rsW9EMwrOs4JASkpzl2JtZojdbm68Yv1IcbfZ29py9zL8c1WeB00aHt5TFHmBXp
j3ib2T68geoDeEBwdhcUZoZsaVolARajLYl+dCX5GylKjIBPFbfs1fYlkLE2nl3+
K4sT2zMdS9nR2r6xoajCi6PFxK27NL5sJhB5++xWxegeVFLky4XRxVpkbvhsVDy/
uPNevR5RHDySDuxtIz/uGXo0tyOBLAbUbWUPcd9UdADLmI+4RtyNCV2PB3wc7VdN
GJDc2dA6XEntDxLO3bukr8lWQ5IBofoRXD2OQFtQjCKC7olkEFUDgMb6VBCGw6xw
USJaCiYUHYIadWCeGRxxU924fuDdBYINr+LbvKaBXAH7Fb43OGYMIHoxN1kpnPet
qICEkWpALyre8A1a9863EOtkfv5igWFjFDo62eiV1wM3MSq2N07sx8MIuR2rKlm7
JHH1V5wetdp4/njVpjJnjnMKxb4+ajm8WH837EqaerKynzZLk0F43np75qJbS1Is
rNbYXZ/YVBb8kgKL6CvXWbdSjqNrQwewP5QEKJjQMc2uBiC7vGCUKme9P7E4cOba
LLGqz+FT1lRmXknQnZyZzMdGNFjno9zqlyU88rhJgzxcnkTcDEOJ/i54aX4Cdnrs
ZBkSQiCISKU/Y2lGwMOMpJZGQjQyPbTU1R0rPwpRcD+a+WPr9nXtb9WKHHsOp5cG
sz0h8/tDV1gVXgtX3SVbGPmgkkcEY4RKDM9Tzp1Q5knCRZI6OiW5AJ2W8q4Ghj1W
a4kpoNsjAkLL93c66Gz91dj7gZ0eHEpVUeaYESs0243UKDIoQBGNDcc1vKqOYUAQ
QIIb6KmtslEyp0NxLq1oj2mm8K5hw3nVa6L8PUTFTkE92jGEIyyXqSRGWagrWRDA
gIqEsgveh6ad5wOvHIig7NmVqJSi5BPaq6EcHEOKdySnYrOI7qMq4BJn8gaKAT0V
1whOh+9sINPqqLKZi3wjZk6bhPf/JKwP/rvLfrluAzpPcBf0QgvuSnbQAjfbLOQr
94X5kbnfSgcSLLc3SeO/hexpRcTl8fsTsqLvKJMEf2mebXwX+tabU3LjM3+aBkcz
I1+EkhG/fPnBxM24YCP+dGj+CoprcsjKeRW+8gpEXvzNpD9OB31phlyCSbnd74A9
M4mkPdwwXR088xs/7FMpz1+9Ix0WLvG4lbMFZVQ9r/tkGI1pMeeYas3cXRi6O9iP
eAB8oY9QOdjMLJU5RW5QtR8yI1RrRhyT+Q80BsKmnvYOYQ42i/+KN7Sn27ry4LqE
7INqw0jfTUFrivwrSoM9p/D2KhrelqW8iwQPGs7NKuxx6/rZUuRF/OdDePVb0T7s
XxOVNKOxgn00cdpTNqspC688u+IVFk7dCPwii/kE/qr/Z8G2OrgwE705ul2O3OEF
cvdu1hlCZWH4sT27dRzyYizpvQErnRZr3501d9xzRG89E/wSTzcpfkXCGZ0ixu5j
YSoOIbfp4HOATeMrI/j5i7cPG7S9llrQ+JmxZW9nu00LQvnXbzZbtg41ZgVHaAIo
WWH/nFVVibqyR/YTfmkEg4WgZKbLkz0LFEtO3Vgi/u43DQY5Mzmj3ANozPhw1N0f
exjAAUOquiq4z+gzZkJXKAXULAGk21yx3RyF8+jKJanZI9UrjTTsPySwxjWbdePD
clEFM+3G2TBQy8FzeFDdK1qwNOMyRoi5RxBstRXqn+3oAHSWsGcWgQINhjHLM4x7
DQasZ5A7JisL+Cdc3aUMDw++DRasVk8H5fFUBl4ZVxchLHl7Q7KWLm7iF09kJcED
A5ItzpLuVue0bEYoaabZITNLbxhA4wi9RdP4vCSLPLLko5cfhLYyIupixbtlQrM4
xp0qLbcGKRv8+KIioIfM2QFoAwcBk4OrUTRXxXz1O/CbR9IlZz3u0ilb/4qVoDR2
2hIG169H5OX1cgOmMpBvegxRJF9dUZoCwhmr8GorAdJyPTAAktpIaDuCC1+uIuP4
Kgtqu5OVz/+rCGW3/Tssi29m9cxFzNM1FOh9F5IqUVg1e3uDpsY2ITcRnu9j2wYo
wtnqFp+v3tYyqgS5YpAtnbTDdXs7En3YnFPfIfmE1JcS96RQ1FsreddeQo9nDDvT
pR0+ucvnJh5Fj9QEyQnYePVEp+U8jzaOfcEE1vMJ4ofN9xyWMV2bDcvkZwNjavVB
QliXaoA03Avbwutb3mt2S0ZcOEv1mAcSF+YICsXQ3GdACdp8K5FQbqUw+gLDzQgc
KWiGgm0KNWdw3lS9QaPg08juf0mG2WEXxZcxCgwBBGI5ZxLWlcgaCrtn56zfWpOm
fOSyT64rSKn0Vm7l1aVcFGDeki0UeMliUlYoKmvTiNV7jjWPBqGC+yhbNJWkcj6P
lXZto2Qn8istqB6Sn3yUvBQ/XbW9FwIBcYqAzCrhuhsssgdiTCNJoI0xnxqauaWe
gCjWB2PDSapaSut+6sNvDowKF4nJYgsDWlkRwZqgOOS+xpttYEE5XHfVwQKztZI/
FoeD4BUo3Q5F9rZ4EV0amPRP544FuWhYIu+SEZyoyqQAHJ54aneck76gxK64yhXF
VPc2xz1e3BXJGpdjPsA6M8Gx0xTJHXKIBG6eY4U//j9OHnXSWCp0x6cCUSAsh7Lv
o7Db+HPetscMKmzzctIlN4URxs1Nw/ErwqmGDZvVfSdiFAIz5Y4o4vspyr9BSxDN
52pCdhZJ/21T22LCrbMZDmBqIbMmJLUB0f3C/EDHnEfj77My8Edhuhho1FlMAwS1
+3Rp1NGtDH5miEWFntxFX1s6/aE8YTa/3mS9ChXbsVf1J5+9IWMwPigSgKt8oUr8
/G3Ds6zb9d/j5T9ITufk9ThUB4jzwyOJz0rYhYMFXS8HkHILKps5NAZY6j9arXZ1
HTLY5159rRNtjkgS7w0MDLiq0XSJBhwy+i3FlRhZgNZZiAwsUtsBBcTdsBL4CSPV
mtls7tH/bY6MU93hbKrOHyYz4z+GAZB7Ne9Uwj1nHPrE97Fs3EcAl4+7T3NWey+A
f80js6fbB6RF5rzOTJ3MCLSTkL5rVwioecXALK5tjDu+ztPDFcS7xZPGMPoDzOVl
c3jPvPjDmahSU1pSAhoKvjhVaUDaijhP3ZDHj/bjROzHAeKfO6lddhCYISwR/qEe
Md7gJfA91HHq1s/Z/U4pFVDKdyyZUW/V9efLbHiYs7PdIF/ib7DmS1HPU8x4b5ec
7YGeBvlx0fCOGiEHH7FGrnf7xHmfKOYcUTeVJJZnN4h57GC9KrynJ79eKwP3FQnm
lX7BnpZQmtH6OGVekcAJH/ys4OYlTnbeOa3kXLpF6Htw86OU7LAJlk7yk6rxJZ61
YOjwD7WnfiSB5twJIrX/lc+KEHQRRDsd7sJlCTXFjAwfDtSKnopNatdJn5hZUUCo
vO1vUAIuROKRncu0WZscPPs5gkNkFxlEKeEaZ1vrOqOrSOXsiUSSK8achYaIOo+2
HWJcxR/VZvw0KX1f2STMY072+KLo1mLhiM6H6KqCT6fQ0Roj4RPTRQzA+0lOcUkt
iP/GlMaXUyUUOLbm3uu+bZVpkqbOodAu5xpxJMYDTVsxUlLCUkJ8kQuiPZT2gdYV
jtI0VyYn5Ks7xBeYJwhZoECVW9U/4JXbSz/Jq2L57KQHHJucZj38qnPUB8fgn6SB
L8JWNO5j6hjc1Betlczd2ourC4xeWoFUVzuFmM8+mSiehhv0qE3QdwOvrZDnKEm9
LnpydCJct08xIzBZ5/KiK79H4hg08QNaeS9Lh6RI1hbyYFEp+xvHsqR37kvOQk8p
s1F7lfciji+8PbZCwr1BLb7988ur8flkPTkbEw4XoqmqGvIY7O4tcE8cnoI0fJCS
ifFDxrKUneYrLqsUCOynPhH/+u6PSZ535aaBmSFObpCKnwYuKfn/JS1Hh+aIMDT5
TS6+0MIEcHK/21KoeG+0GCGf5gbjak0vxDvrpN6M0YTrauUjdjFYJ+XhRFn7bgfz
XaAXr+tZBm9ifnaKwrCdF0PyC5tPIV4gIu0E13SVFY2kBSQ3KuMq3dEYqpKGBe0F
emXk++dwX4np94aobq7rsNno7jju4WGa8P+pVhWhxQeC/+8lFeETC7DWy71mUKtV
xsbkjFb/zjJtXIsVsVDk5rcLW2AyrV2yhXPQgeNlaaemdcJQjlS137ncAF+u0psJ
EIrkOlfdgYohVJNVHbL9PhSLpYiFEnWknnz+w+2R9GTLpendNKwS/kzbHS3HCurV
bT1iboYZ/Puy92tG0oRky2B9cqsIYKHV+kibsN3DcIs3LFWowMJZ3PIXEZKcK+6k
aF/2bmqEPBQb5aeB7bVb4nJbfaCWiaXCOhqwjwUATT1QRj/RnkMcAOB1pzItmKok
GBfMp58NcqgGRw4f+UwjC4e6JV+jbDrFGxS7FcKKPuhch19vYnYD/EZHgUMPAV4G
uKcCVzTSaFD8M9VXtmTfwStm1bSQxc6CzSeH0ECPw+Th4S8NKRkNsuwLT2larggA
8Sn2VA5D0XfHn7ApzNPj78iHqWaZFCdXzVmHt0JkG5MN5xBQVdnAnY/H5pYB2E3P
r+1wl1g7NKPlqT2YFZYMrlB2ck7FQf5ddRxpHfQTFx/X3M2oDIadQdmfZJZujJub
Fs/ZDwfr6i/HsRzl1BUDYal2IhwQfG5JPADl9K1f7znc9d22vLE5OVZsUG5kkorI
l7RQPZ7TWE4SLBQpqcZJ+rTsW3yAmxLrsc4oeVViSA+er+V4hTL8YZzR2P/v2xJm
5hlBtAf54jrbB4m1jqZ/a/ZnehNnNZU0GuoKgo9aLkZh8jcjSpIfdvq3JwJgOrO3
UiX+YmZxz58/7eCmLquv6YcfbSM9xrHvVRdTk4dZTtGuQfyRRSgS0qU6vfKVVJa3
wrdyMWeQtpXf7IbroWTdxtlHs60NH5qdrqyBH+llgzaEvM/ZJmKKYkOoEQ2VEKPb
HT8Tug8K4FYkt/B4JC1dmE0CZQUWNaLS8jdAqxLFKrtV145DP4XSfnkWhdcLMb2c
xzPX26iGDCqqLrYY4idAzfholInH/sMMycE4UjG4S5qNealAYf7cyigsMtBXlxPc
+x6+Q711Ke5uYaGE8qu0F5H0e9/6+BDXcbmtB1MS4gqf7t14rwO2dHBNnynvS4rW
s9pTvlQxyzzqaoQaWgYNmRBt7wGbIfEa/wA7ygI37P2oNTfU5/TeHHEpAv5hq747
yHUP8MGi4oR4DwGg5GoT3UV7NNlprRymyUC29e6mx3aPHh+PWGPNhrLFvSghKBZv
kupOnIXjYuK0O7fwGGfDQLwCwEtIxwqUBKypy0icqpBdffpiz297LPd0KFa+CvVp
Q9i6CnmLjLgSd+XTFEF8HJ4AvM5vKlRp0n4pq4qBN5nR5tkxBNEHbVMnocgrIncr
5rMGzzAlYrG/fkjUr7CHhE3OtA3IBrO8n9Hc/A6x/G6G67qAHcEseSZoA94AyOOr
ThU0vwgghgbCphU8htPJcJ2OGKx07tZxH+ckowXvZJvght38tXMPXtoucj7ZvjQa
u1fWXksr28J/dHdOaXKwB36KFXgD1zpUnDN0wk7p00mw34ZYuFcqkU8e3HbHvBSI
y8ebdw7LAZjCK3iD/jsT/3nhOBRa/T1BN0yg+D/lu619e6Q0/JaD1eatHfFCliaX
uLlsxfbJNLzHf2XAAIx4/9qHtAeA7MVGSB6GooIqSC3Ild/xiq611i6tLnVEw0nE
ETy2FhFDiXxP29gA6XN6f+qr9Z278LWyUa/gk5ugLUv7DCpOL2Qi1CYU3iqdg4ao
0V7gjVGoIevLza6AdhNoTcCWGEYqrT+1fojfhsbJu37VU8f/2x1R/7GkPhomaWML
w8iVZY9JRfu5vV+Gz6fRsf97cN7pwL4tnNcg1REpvkPm3pUWyTodcp4JJtcJ/c8u
BLNBHsKLTxSmVyHHC8tB5ZLnC2R6wA6RFJl6tVYMyn4pjNUgazag7a2LK/NyaxWM
doVeH3CGsCSyy9I/Lh0tyyVjs+WgfePMstiaIVYNjGJPymsQUdU2X2GHWOxv7xja
vs9n+HEVNbU0p5khI0xYPJXAFsi4CRbnls6L3PIrwLajTHLG7zRIBUiAedRxeBFn
Hb4MJ3DjOUftHqOpYrlTVA272ioen/a8+XzaXIE4RspLkpS9bRgHlJv1BQ5Kyygc
idZpf779jseHpMJbPEF2i6nkasBJt6bqiNWhQ0ax6KhqZIVfzlNc7CPENZctrw8O
CntWSpKwPJayN36mT2dq6T1U0sD+vTcBvXIoMMTvIDpaoYQZQicGcVIHp1MNC3MI
UD9KmvV6BmzZUWTKe73oRQnGJMoDyzU8yWTxlJcVgSwmdZpb+99iXNKA7At74+Xr
r+pDyd7m8ha8pV4xChllCgfXVU+VNFMGt8khT6kC0figaivSdtWdAi4nHGNazp7D
yDSd7nUXwUtofNx3wbELeUz5/0Krgn+ln/VMfMTss1WbLBB3+Xh9q6EmAf+Q2Mnj
NWwytycE7dGyiFiDNTRLaHqhV36q53ct1Qi0LLeqMusB0TYKR0qKRrg5hPNkp6kq
Kwcw9YMyb/fPeMdBYrFJ1I+g4f8BLG3YEm8yTzaEB0SVaGgybPnq2UxCcORE1UDV
VJT1CvYUj/WGkn3jfW8wk4HlS6uIe9bFL5LxvkTnyQvUydnPHMJWOjYSBMFwSMLw
hGtx7zKCmNRHegDBhdqUGPN+ZSQ5W02WObzQnaJmD3MWRbJduEldww9Jz9CC/AMK
19H0REWKPGwDLB3ZoadeNDOnYx+qCSSdvWSfb5qIMlvyEB8HNWMtoMUnE9k/WUMh
522S/tXhjas9p3d/ZEChlfh2cdGL+88gHOzMEK3OlqEOtaPsoylSyqtkimYy30Py
76nKPDubzLUAxQYEZtzWx6ZaUmrz0Gu4KM2u4xMW7Oq4AG+60In8Oi2h4JMak4XE
hELasyiwzHQYPPeCPAOX5EbRCWC1GOr3HrZ8rayiG6jhRCcJXg2bUXSw5LzXjlT7
45UuaOj06yrvF3FQnj0dbsJ80AnC+jtRS8oIP5RePOWN9udWK4BR11rDvyJQeTs2
E1HVET/iP7bL9VHxJS37C2wlmHTnXEtTKPJJMLWprT8kwWc653u4o0mlGGcz4Vi7
Ky9cQX8kDLipVqTW+kfqa4eRlgAKTU3gxTQuxgd+1EyJeaVj9Rt9krBQ9hS/HCuO
RKz+OYFFRiwwiRW2/FSW+Lpkz2Kbe99+ARDCiYw6kkzQEG8n5n73dT1682fVgR+B
6QltSkp8vzpReR4wglnVQdE+dtgGozW8jRSCXzdtIagrsARHp6JiuGr+idBSgjDv
UBa2O3BfFEySIIxeeGaaBObwBIZVr3seeQ3gNvcmIssZhzSW3lVuIaBP9k3oz5E8
23Ux/UbTplXvsHMKkeEh4TtOQYYLn1t7fqdYeS6rjnZ6PzampbkFBIixfNWtrBVh
YbPC+VZCELQX+NAG8iXw9QrwP5sZblrvUhkkdcLc1wN7uXyYivlLTR86Y59JcTr4
/cZ9Q+kiunQkLYn3CndeMvXt4xkOppGXANECgrogo+HLjknq+NxdbLFYYawgk4T4
t7Gm6wIRCzdpEAM6Aq0T7dAcoTrsNnaeaXevpuKSpvgPRR36kYhy7IfNl0tK+nmz
FA2L6qVE4p5zRmyWLCuUzbpVxXvTmoB6xonlAqhu40lX/YauVq2rOoiocDFWLT5c
92gBfWEz7UffGGLnSNrrWr7wJjE57SLzpq1i0CbDpyQV90boqQWCaw8IG4Sa0wKt
ITsCI4+N9khbLo9SxWDtj5AkTGPMntNa//XsoJTNbLkoJdLGVhZUAYdG3mAPfkXP
46aIFmRMRmUUjjk31sCN/++LDB2vYe6duINuWS40G1DKzfx71eaekdS488vVF64G
J/6mnxi8IKCwIfKNvUrKqp1CuwzVZaT52yGuJIWYPcU2s3iFc/QDEN5t3qyEnJ1J
kjM0eF79aX7hy4grxJF+OaC793H1n8+ujfFo9UrQZaBUQrTlBNJxYYaEMcWvIfEZ
PSBy73JBhWHqyBrI6kdhiUAUOKgVifv54ByKEGnYUIc9kesOkPHycefCh4c1mWPm
cLoubF2mnCoIoIDrwEvA/Dz1XR0zeYWUrl3RxpJgIceoAMnQMvT5vZY+I6FLGg4q
hB26P2bDTvBA3Xp95Cd0LPJyjawRSC4zSOJi8NrgNgJDbtQ2LJhPXWZaG0ukC0CT
8X7Eqtlyx6nXz+omMT/c72K+8NyhaT5skGvW/wRm1zOweqFaaXWz7ZKON4wOzIRR
9r35rr11CLc0NJ4RF5tujFUk6alNZJF+75kTt7VoB+t5pacFEodszotK3ePQq3Hx
9EZtTAIwbAJVRM+f4fYZdVJIVnUfM3lJY+0O6yC6VpzrWnGCoomMA1YQtMFztRoX
jdzjXnudu2QgyHTZzyVTpWJbKE7fzTMIgqbpU4IkxeQ1+wYHasUI6mYj/mkxpl6d
rZxb0nAJXqeGSQ/JvbG6ikX0dURCCeudOd+dfVF6fWIFgxomk+iMUyMQ70h23io4
6A2unjwyxXNUMxcesxGvFJgwxLKrTqP1A8awhZEShsEOsYK23Q1v2KuE3EFouJPK
CgPxqD2XRsP/CVKEqT1jecaueAjBOoZKDpHB1e5R76J/mZQHR2xcurtlNGiJxh0V
TkJEr2oKbshlC6XZaQZFX8cFRoz+vvxUOL1XanJAjwVh3TiGoGi4F136aqe0JYRO
T8EriFQw3fKmXHOuU7gsRta1p45+fST+29/3h14saJ9XHrkAIVamQTOMYUQ3YC8o
XZWv/BMesgPHLprVkaVqVIgkKVgE8YfC2NAcmAxD+YoHjjbCkaGFBq18kn5ab8ga
PI7qFxjl7eBxESVJ96Wft5lQxh+/x0sP6UuT+Xi1o7JwnCzOiX7ArtAH4+ccvCs7
keXBusytVnnTPWxN61O0sgEMGBrikKLftilCJ4qdyagLuZmxItLtQv8JkRjM6DrH
dhHviLRLPXccR1jk2kVvg90ZNmYuGKJ1OZ+5DMPnbcnqmbgRmwNoFMl9X7FwWu95
XGgBGMN0j+grb64Tykj8RMw78zDKwHCm4NLIGWk2bzEapigYQHCB14e1JFUwT9MR
826GIys6dMOZ4qL/yFblLGyNeuL4BmfI0icb15aiWr1Y1cOWnNTMVWklUJr6yqPZ
xBYNS6X8K8fOu/W8yq+6oElB49TAvlFibrjXwmtLGJ+BmWN7qJQ8qfbvph0+xjcK
ruVRcF/k9fEt/l/JJy3euu+gnHR4wdRR7xXV/gV9ZYiHFB+lKSR1Dws9EPD566qv
xE98wMrj2nJKbX0oYBlMvxOgjSAyDdJZ5rwxsjux8+2vz2/ppfyKb2aADDeWreCU
I+eREwhStyHEyCrY1yinXyIMDLVmz62KN9B6EkBpSR7vOtkrY+vhSKX6fZhRw9Gn
adWRHPhIKC4XjOrLIofdVcCgxdRmEZhKB4xp8fSJ29HVCiIDXhXS9Vaw+qs11RaB
7M4ClXQ24QhZj4O541hYkuPJJpL6ZprU6YblVsBfAAPRbSxYuD858BjGfxsNcTw3
sOl0gDLqBsNPhUFWSbJxy9XRlZdA2nOg42/5IgsVUQv6ds/XtGu2UFQGqnFODzx7
7QEBDp6Kj/6BQBoD3Zoug/s9ORhkLeQDIekNv8sjme5JJ9TQt1bTT9YJrgk/gwTT
lR0WK/cOq5BU3KwVhRZWTycKeW+FuwZ3FL7mqL7CGdRHw9nUt3hx08jc3gUBvUFb
lbgsyvFcP2vWPSvQB0o7Y4etWVdPEzVWFwbNyS2t7bwvnJX/L6h12VUyV2HIlxkv
wTMKoIziTT1TiXeqoCUWZhmvgcqy+psEI4n8dy7SU7KHYR2NGzLIoHC+Syt5VyXf
E5NeEYy3n1CPSWGT5ev/xQAxD1vnxfzDijqAEIskEM3V2MvRuVNvWwYaTTuNz2GL
1oyPughoGhsogJeEa935mnirOnEq3/a9/Xr8c8t4njHOwN5HnlthZx2BUxE1bCBq
XXJ45SBQtO1vBTjkEu+6XdPYrelxKow5cxkKD/EeUpb0EDJLpsw+3XxSfAaLQugs
0yUrU9ikdoyzDb2iJUS74jmCGANIxWgRda+cKDO5OFDITrZinMjupRbiuBC1BvMN
NlsOMfEO7/ywDuskEq0KfyWGG93S03PSQNjUGQ5wJPf2b6UZNCUaoppqYLM0kim8
YuwVnrUfiUKIWkpWb0baImXlN07eX45uwsZUiasrgwpZMgFUX0+qzdGzm61ZIK18
3kN6c1L49Fq8EQGR0pGI8Sqi9pAeYCPHWdahxuUXXRUJcjqhtPIj9VQp8C7VrwuU
Prp5H80NLqfD6ljSiVHvo7cZ94rtZseOdnfetnXmpSpbeQLmcu++AofPjnU1HEND
K3D/98oINdXvPB592NmZoFzls90QuLpDItHzhQC4LoA6yHKtelcpR3wVJ9pbNVJw
bEsVKaBm6lUZTtivY5H1fO8WRZg8zbVE6akaF8P49hoQjuOLiPfPaUD17/DEVFWM
7QcDSiQ+PqNC7KNH8WqsqfSL9x1Wro2/rWwGpff/xivLm1CS0/VwchwDcAB+vf+0
IH+Nmnt22QQuJlbz5Zmb0QB401dgjBaiN0SOj3IFw4vMI0bZOSbrCl1+HYSttiuP
yntQD0kVAnVglJU7JFpkE6xpWOZwa6y8QtSC6Cf83yznSKO5l8nrVCSeq3oF867n
eQ1WPmL9fO20WB1U6oJ0SsJG/QJozTlswsCUNhekCUaW06/5bq0Dt1mYkBgZ9MLX
h72hdUPyi1z6f4bZwX8QJ/KvycWF2OZeQJLhMIFtHAtGze3DO0XarLcp6xOyImXM
/UKfgdnfVycjkyocALPPDKteyt5A+R82RVpIoguj20TwIV2RxJxFXqUkhWyR4/Eg
PJqMzhHvXEQmwcr13M1V5vGNxuSTvVthIF1p8tGC17kCqhfFoaGrjsq4hbAg11RN
KV/hj+AZaVWHbTpTIXZeI2SdUzJ6ZefbK0oHyVqX+pm5hSlqB+dZDcYOTaTTKopY
7Kq0ZJmlXJsjjoPk0YYYNkX/3WSaXfud8QeNd12zOzyzCaOl7fPnceLY+tvcV/cB
5nWwjmmDF02PR73AS91WPN9v95f3m+ykiJaw/IFO+UGhx20UJcK8OsSKknWtegly
k7XPIqBUmeN/gW+V85EMHwlozaq3q8vxJ31DvBu45mdZulopwG/DgPF0S7vGGSCK
8RLbJADT+LTR7C3pFy1oAeywlbpVJfONJF9dSpAfc/x/ZpLDRI3Uq2rS5OKd4S9Z
+/Ve537ZOmsGECHg7leozZtLRpT5LQpraCEWAFDMLC9Hudaz40mvJmfc1DyVq8Ma
g5A+hwvTYLmZuVXxjlB14ctc+SoEFrYsPYszYlO61+hzG+tgahS9+FdOpNZUlqrN
GKKE5Sg8wnRURGRKbwMRoKKaQgyERbLq38601GeoNQkIieYjVEBq1sg9ukX8Bz2g
oISAJnW1fYeHTXhAzGANx5aoB98UteL7p4vHuJIOC7loLtPgX6bMC56+5QJ+Ly4d
b5Gm4ek+my6cv5/GQmNnSGcihy40i2/3nhDitsthjs6Vo9uxywZ1BI5xTi2E74fi
5v3ApqlSdlV2X/+VBrN2kh8XD41FT4/hkT63/PQkMQ/utdRUiSYDQU4iywp8P3XN
TgzdI1yI7ymaj6zZzejXcBZ2LBdXDjP7lpGk1/lcXDuyaQwVjeFxgf/FFC+4vB3e
69BdZQpNm1C3qp/z2N48OJxWu4fvAwA1NF8wlvBNJL6Aqvylj9dMA81+bSMUVATf
WUV6+fYOSyEuzKkjkvzSwX3WyLlbp+q/roH8vZOSku61OTHrS6h9tUlcgMmqwpMd
PxbvrmPt8yb7hsL1jXV8bnL6qcEjuOiLpb38bjZbW9lYyOtl4Tq7d5O2dL3pQj9E
oWy+mrjkvDz6lDER7D/d6HL2gr1eyqsuoFdE9rCdWeDEXCeQi5ahJcE7GkevOIEw
J+DnwekIjeF7RcH32CdPYdp9NioLzAS8Enaj+gX0WunXP/m+WHKytjj7dB8KNS5X
nU5hbNhr5W1QAXsbO1+fUDZoX2BxyfRGqHYMVNbWW1v2lMAexR3udwMSkhMszPkR
9STibZ/+NPEni6NyvOwFEK4bR9hGXTS0EP28coo4axTCGREiMoHGlBUHrMmRq/pg
Bc7QX8MdRK14tCK92G//MtdJd/lniXz323ayfUYOAwxUdWJ+bdDrCHQfOQe9/W5w
hHvOo2IYo4fA3a8LHphawzyBLbXwHkQ7awODHjyDmAmprI8wcaKpjhVWplfunQ1y
lp77gLFxxvhSDO7kc3wYRkV1PsTbaMQkDV02NVACrMP1bXO0Pg5CqljE5wrlOsdC
/u9EnlOXwedzLgHFYhw2yEX9dNiBRWx4iAWMMrEreagXYksQBJPQ0c7c8hhaHsIJ
i+/o6EzC+Ik/2AGWuCQZAa+yN3T0vqVTA4vx8QUX2QxTAi/i1a2A6hybI3YSu6n6
IBtZE1icbyo/B/VVzbqsw0Kt+otsWyXjBB+Z0xj4aYNtUotzfg2VDd1HjLo82ETy
8MCtUJUvtghN4ACgNJz6w4Mxq8fYnE2YU877IEaB5TW7fBLtJqpY78IQD0bG1nsS
2Z+mcct1ZEDEhhuvV7FiwkS3ehVzcHSi918FzIQjv3im2v89NE5v6G5pltTo0SXG
mtN+UHKYtH4gPIFpCuV26oKgblshIkei2+H2jR35sRbxwu/44aUGleHyCXYc4gyA
B9JL5nIWILcmxPl/kSjc7/VP/Y1KNaJJA9JWuF+enE7O6wvEvO3yOYeAV3hVXn2U
4mkObtG5ndKU+aUkdFYAnFzmBBh2g/Ql3D8vIjNkMwmTgpdLRc8PiSMOUjqJ9enD
j6X/qqpRuGj9SizyF8XFVDB/dUVEAL+nO1EEpdTZf3EVHu06HefzqCaia02ia4Q+
vva82rHC7BsKoJN3P0Tyvy3/GhBCD7G50/ADbMIZe73hr9aY1uL2WnleTqo7usXe
l2XcIe84toteyT7kxajpTWsv07jxYo1xrn7m/A6KL6MgqUgy3V6hW3mXlEqah8PZ
WOFGBbwryJuiSA/vQl3FYL1UPniWjhmgQU4QbfGw+AZzMyxk2rJoCKqa2FusNPbx
qmh3sTS3V5QCZ16MmUFQvLowGCQtyUTh+suFV5ziS+hltD3HsYa3w7dH+l0caO/y
kipRfGe4zXDD7oS02NY4LoUBtZcvloo6f2cSVS5QKJ28UsX5A+7hKDJJCyhlcd7e
A9n8oYXxGRzavAfmaLCOZU2RRjSbfsNiXyaDGtF2IixpwFbvnBgHqWFdC5PM8y0G
e+J3Jvfs6txnJX8PPXyDvWTeoECkAQvVdwN2sHaxxF2JFQYGdyHoKLJORjERh8Ky
760CWpji21ydNBQ+EW7sktdvgVFwTuW9wkdYyZHVX+4KnDIn+o08hoM65rhSL5Tu
/+WYl222FWRGMgs2pI//tJlAVo8VrGbF0URiqW8iuM0MCsiiJLN5h2ZBQ5ebxPK7
un/PcFoJ3c82nnjLO8ZUSGcK7grvPzqP7I92XZbv/YtZn2KTugKBy5/jHamAJDIm
uVMfUPX+F1v+ly6ZUFprf3i1U9BwLK66GC+tPrN/NBHGmiATHZ1Ltn9FZPQ+FrY1
HmT5Iel/9tkw4iw0PYoVRXX9+UHVINTZB5fBukCpSij7aHZOTivU0GzayCuYgM77
AyuoYBN9d111xnJUE8nZJUrGoWKZ52xm9HT2gJEON8QaOUa1d1SgFWq8x9C8B/8b
4Rea2/Jb75c5yhSfrrx7/BElp1t/Gq1gwvMdIgVM8CqCZjIEaLndrp+IWMj51m+H
YtsZ7NkRfUu3KwHrVD0+rT9YpISv7pWDRgdjgGhb7EL1Kv8DpAFw0yES3mlLGuV+
JJeVZUSoKzoMNPIU01Ile28IJR27bXdQ8DXioz/Sl4S/p+78lnKHXUpniPfoJHTg
LdzMbGRre03mMTNPWDFH2g58nOYYtmrq355+nasgScHNrGBdWayH8vqB+V0dGOHQ
a+gfsk8SjZPmPOmWHDU/A/r7hNupGlhk2DxZFqyDwHnbaOWwU2XTJ/rsq7G06AYR
AOfKtLbgmxMBrRVauujehx6NVJ/183CSgtiz70nP76o1jiP9j0AYOu7MTHVDDP0n
C1iiAHyEXAYlzVTfom3YCNFUkSae0dapjNJx+eefIvhADXguZPMuig82mRVo1LBX
9rjBWAL1I0abmTih926tkpof0+dWC/cyul/rmotf7rq86udYLN+dkqhoRrhkmg0v
Zja4HDHtaboMsbgnzXd3zisDZublh5wcTuvIGrWhISHkLKh0NdpiyxC8jF0LqlKE
369gSCmoFfTOA7fcNWwIHA8R+ZDZGIzwiZddY2XfYfqQBnOmxkM//SqNMq9I2OxA
qArcgWBUm6wVZyknl2GJFr8VJkdeHQ/hvZyYGOJRx0ed7hwbQPhPtPlabRUewVbB
GBn4mbYzTCHSBT+5T3LU4vig+7+8PcbQ26WbZd8UB8mg9C9Ls6jl+zSvRS6Q6hSU
BvGaqTlhguBaKRKr3/EX/RU53/BY3m7OUMffhtN35DZfESOyBTEaL8tQcIyAqHv/
gD9kpi7BkjQnJW7stbmeKQ+vxZMj7bUPv3GcdMbgy6BPtaO3O6A0VPVzt6S3EBpk
vOID4ROQaP/+LCQbtcIhC2IOnw5YLYKVhDgOSE7pDeKepYP2fWCabKWK5HZ+lo/M
AeSenRFoA9yVJsb87IOj7QbU80bGzyAe2Ef4shbhZ58+b+L8oAUhhGvBb6mIl3MX
k7iVax2DhBEp9bIRlTirqyaf6xw855WNwBwUlmF3oT6f9HarjwljfzolRzfiiG5h
sKuEip4B86OftFzBI9gm510MPfD+E9ApBRjh560JU8JzvOsrYHm6r1P/qCxLnhGs
IQzpnoLHY7uBQRKrSqrfP30OM5l5dTVlQLTIPfee0A+og+1zQV+UvbtM3+OlNVEe
lGtcJ4ZcPnazt72RFMElEVPxi7C2cWe4cpk4/zUdW9kygCDQE/NjEUTpGRJImzov
yGWX3wh/BSWGykKvrNQpl9G4Ugm9IMq6lvhbhCZmDK+qMuaTS3MivBmHvG3IyEg2
FXimOicAsF4vnWZUGWYkR5eSEQZmb115Lk6SLd7NELNM+Lff+OGVsnbEfkXFziL7
Hraz6GgHGpCxZDbNlOefDUt9uYCxt7vwXhdB+MUIvy0FBLOAsLWHeMLmueb2/8kz
hULy7WSS0uJrWjuLkvV1+sCxUPk/HUNVojoIsUQotwWcqZeZSTBM62YzR1BLPR7b
u6a3TRxbldPXS9Jhdl0NkXz//UpF18j7SARtMu7kdJqLONnb2vbqyj2UjybbGAxO
oxd9Rto9z8+iTXGDNksI0kbd4dhEtEh7g80iWR3BT8/saS0Hcvk3TpQl/Oehqgv2
Q0o24LtCMmY0DLmT9ocd8eN291xJThZ5e4N3lRe4kpmdLXXUSyTcHiSqKi8M8gJI
5Cq/wudsFs8U4Uev5SJ+aZOn2SkX94/NGuZBkLGhUPQOAnisoKRWp2Qw+Tajk13E
x+5ADOuWYovga1Yjf5a1CXQ8vS0DfyekFxL+f8cGEXkEdnMX1fsPUNkJO68BG9AF
9qqdPuwBc0PNtgGcCoAdz5NZNijq4cwNvdcQm5T72LhQMpPp7Q+huXQrnY/2iHCG
tuEVZ/+1vL9iI4k//Eupb/MubNW2J5jU0MZ658xmaW9e4IHxTD9uN8EEpxC3lxeg
b8HNqJ7Sxny0btTZa0MMqP0UQ1rY4P9pZYhSxqoQFg9uCAHBLBsJo1HvcVCTBAEf
2XLCzbhjB1tXE/td6b4RTJ+OpbMY5BUbdafsKIayuYSzjCc9bf8UVp+IubvJay/H
68Rc62hWeD+QNeMajtd0KTGAW18M/jdo23nel0tu2bwLWEFC+PCTwXfrnrk0YcID
gzg9fsOIKBbiEXXQjj+biNw35JDdjJIMVsV7khJ14K0R6J/9lzsbUwJ8puhxI7cA
1wu8LtNlNgebRQwj6K02MlBsDnaFIZOiCP1pDHYqpYNMZkUIDS3f7rMQ35AjYqGD
UN67lWSLgDdHjndSgaPmbmC0PooX141X6TyYKx6RoWNlqohFppKAUv9zRULL5xqh
QOxqZ6Y8OV7Wv7ewxvwRVJ2a4coy2rvLutBIfQIjEqwDRNplbJcUH4jhu/W/dzVT
Ni122JHIEjjZtZEKHjO1d1AychJACYyxqzNXp1JIc1GkWZ83mbkjZt/JK3SGYayX
qCenE1P5rusZX50z864QTGzJckHRR2D8Xv1Dc69iHTc+R4Ia5jOI1Zs+L+/zksGF
7lyKXtmRK20wFTedjy2nP3YPk33COHfCs+11TTfYQDFc06ihWGiN7lzbpKa4GuSB
NznlSfzwHyOcqQoNJd2xFxVDo+dXNqpGSE8Teo7hA7bZC5IU11yE+lymarAXQMNX
PRVGlESyvmRnAOT1fn1SkpK30bLQsdxhYtAKJ1CYelmQu6MjGSPYTJMWoph/Nny3
jqrsG/UKJ12DTghtd60XHGZKzCHENQxgR5VxuQjGY6Fn4yOQaL63kFm7DENNkCWj
6lNVGeLFJd2Gr4O4SKEFgKZ3U6pV0mRe6K8D2DDTfKxGo+W5smvaK36Btmu++yjE
iPzTfwgLOs85VHSwwCBoAq1xwzbaBbAC5aHoLP7/dTDyqB1BUx88o2K69MtrQs3f
IMGJULyxd+y4luHcSHeSatcEoZ9TmeIntbx6TP3pGPYitdbzT90AA6wMXb8sOxlJ
HBDSgXS2TitWd9r19fAACVqDYl0bHrhuWo1c5URYjNlVhf5WiJ8IST3uAzmkG8tv
SrNzgPL5MfkZW3phnDxKLRboTH4QxGZiGgthz4kp2NkXiDleQ+KS4yUoZYpgnxUL
12OspywqZuEODeMYHBCPqeh8ZAj1j7Mxebq5YtU+aexPOsGxIavmTM983lJZduUk
N7Pqdf7dqnFWj2Nq7uWOvSXxe14tZ8nNS12EIB9Pq2WUcpEnt6vyPVJYpJAeLPBf
VZjkbBejQSTRC11TuTQTAvZYd416EwnRYts2reBQ8Ogm7ioIAIE8Ga5zYSqpAuXM
4WJNOxGJccePUadXeuRUKtkBDD9gf8kpi5y8FohGeoRd5vx6XqbR6/ScqcdVGis9
LGHRP5vfRpdM/+t8usfK8N+MEbFrT0FNo6Kp/YnKqwYkBmcSr47Be3SPvPXAK3pN
RF6pujy8E5txIW+KsyRPL1TFo8gWwPsP2P9yoONVfBasrxbf6blBZPZ6yDK/eBMr
DRx42U7vPn6rkaa6h6f+lf9JcXi2E4hghVFDA4zPV+7p1OehfEMCc1dHK8Adejxa
X6q7ssUB0x27KV6t7BeXavbD8Ca70ntZ5YBP1U0jUSOYiTsSm2/2Rmh0zvPfk7xS
sW6Fi6Un8H329t8Ghp4C1FVDz2PxRblobmo/WFqXYLC6B3fBwzBCXbBazKDm5Xnh
gDPMLREXOBL4eejW9u7/fX259qB6hK+CUFRL7Q9NMwf2ANN3mwEf+VAIY+vZw/Td
Ek+HNk6nRAqrcFUWWqEYBYY4cGhI6PFDfSu74AQTu+4vzHqicLa+Emx+XfPneXv5
mRVcgvHhGhYLkFTZWEkVKd3l5QJ9cvx9LjnVLfr6cdHV2KUaMflgeORQhQanJvWS
lajk6ie5HMqUx9WuxTod2xhE1vfBKIuiftjrVTOCGCnzGjLPSjMbGVY/tKFmi2Io
EY4wp5/OHbCRYbSd8mBrWceF7z9fmdJAV83ruerkHwRAeajDhM+7bUnKUIZefgf0
y5aoxBCsJ7QWxLjy80MVUEQ2ubH7AB7mHX01sbvS1gPgOVF3AkbygbvuPjo7HpsE
vOxMMtVxQ1GDHIV32Vv86OWRI+j66OREHTUEG0HXJAZGK2VrN28/l3U+vzidcNKP
xj4/X9KSlhVeO6PMfdZCb3xte4+4tVYHhmM4u3Wj+wL5LhM90TwVxOt6zcyJy+oM
Qhz76PEufN8+5i7X+ms4lE/XwevaAIVyXTSq2TMUKUVSnzMR51Ix3ayS7h33pT/H
JRbr8TRzdpfbKDJKqUQ0+BSSf+Yzu8rjzScvP2gxJgxqdpG1ZWgyFRkAJwgdM0oj
5pmUb0i9HsiRcxp4qsuT3SJV8DvywY8fYG83nvl/MDLjUUofNyZCgXPdMk5kD3z+
PpivGu9zR8VI19Jc7VoONBC9aQWVLC7XmqjxX4W4ditSjE+pVJZsoKIB5bTpe31O
vg0nk3Njh4XzndC2vXWIlbksl/C5ULQ76Ae7gLIWCmB5EBIyxU9B82FETz/PBJh9
dAEAyw5uoU0Z8yNUWBIBfmi8Eu06Zjv4TlG9sEvbBNDekuniBn6X8svxkZCQoeq3
4uC5tyD/QRVJmqEoH8KuGz3GEnBZWJwYujAF7USZoKltHFdQ+hsMWBaEinFCJjQl
f1nFf1YSKQoc1uUne1owFYWSyttF6p9G9ZLBLe/TkKFbiWkMU82G59BzOwj21Tq1
eUo3AdTYmTFUzTDXcSaIeIZUK+PGaxIxD1zWKvnQmUZo/mC71PjZCJOrBH89mPRc
TI7l3/9i/GEk3JMkJnT804RZUa4MfI77AUVMC2uA+iHXItvApqrGgTGLZAR0U4SN
tCQEnwVr6lohYT7tmjLh1CCijD/kqghFK/SBajhbvx7SNULBSLMAjHzo9cjbUnoA
oxjF4snjodUUlKZiooxuadWnkr7RwBA1QCJTSB45qyrf/ba61DVWGvExCoVHJa6y
sjShuuC88dgk+yZHNJei+aj6DoSODQOV6JtFbzud5oCxOHJMloUaoJzFRNxJUI3j
QGfyWbBkZZo/bOm4K1jaJ3CDegO1O/6R1RBPEsKG+1TwZoOoEPPPytWuhEgFsBRt
Uz7MUIg2SNeLQjEDbtj4o42+OF0MBHHHTzY7AI7NDbtMSVNjW2jfViI8E1yQxVZj
Vb2R5TLeZ/ffZHBx9TYJXg6wiZdj/Rd7/j1t8TJCmYYHwnSPJbHZYOA+s0vQ5AU/
Xafm9Aa+SZmOpZW/GunebjUO/2hesvb67jNF80k+7UuQkNVYpM72y6vPz8oed8EH
qcq5I1Rnnc+6wjeIvMVouvvc6PgRZ4Q0iN/s3uOxCdtQ4ecthmvpehvYNRYrZ1ZA
31jpoJD/j+5woxzy+k9mZRZdmS6TL8Ib+NgpX1RM5LJHL98r4EEAUNQDtpU8lJ4f
9wiFCn5brCOz91Od7ynbeJ7Cfe/x4VipmjbiZN3vNws2vNjtyJtdmPk1Hy9Npezk
6T4FAbYiN4TBNHtOL8o+SyAz08CLahRfu0VM9VM8mB7ZCXGMO3csIEEKz1+5Sc4d
CfmY2r6xUtdVSrpNE6+KKpD4qaYpGPjGTodLshbgH9s2hhFJVXvwhhWYwXDw6iIg
sO0nMNc3U+dwVxCEpekgqRsXxOF5NAmITPb8cod6Ne99Tf+GU00uFIZLJh1jHA47
GN4FqqxHTzfeuJ9X8lTyxgdUFcgQh1/TX5yk+zuqkQsk/lmq1ZchJFd87Ykl7kRc
0sJYdVX92IdesLewhTi4QfzTUrSIeK52mfJVVYa2loyxVLTSrwFf+9G28EsvLePy
nbDZwf2kaF5Y+gjTM61LidzK84U/y0rqKZF2L7ZYt0w5hGT5aXVxkbPcGI4QmAzu
v2wXLor8Xnx+aYK9mKxRhYMQU3qZ/D1OcIihbYfzBBqkJ+Cv3UPr7tu0ebgOpTxd
LJ/g/LH/Lulft4yV1cdpzS92vOmh/NQIVaqHs+Crb+0LwXBw5FZg0Uh3vYVL0quA
LJx3kXRXcsx9pHMq8kCTWCVnqhZbnW2x3j1eLVY3AOPmBLWrNbiIenGsRuJBL6x/
WxfwrEx2Tv7kVdMubq29oNJqKTh6Wz4Jb1jlTJTu22T0Jw+j9NSZ/K/m6/7g8abl
q3xvEE4Tbxwd9Bk5sy0nthGabMSP7cXsA63ZRurmHK1jC8E8P1iPgnW9ms3bCrdB
OeRbhhbDFbbXtt9rYkUQ/b6mTZsMhZ4ZxJq7wLthOllt9U1a6cDrwYcl6rgtSdhf
JVWhSGpzDz9G5RKMh8OHaENxgl0K7lMmKs7UDA8r9A7J81xnKvZJTnhmiPOYlXyv
pGXMePEe3CUkXXu7gF4UWGBYpH2wXPi39NMzjOo7HT47nxnvOp1D4L80GXPhZsKW
G0hz224ZIaVZGDXEZQXmkcxkGe/BGUT6NzoHUF0xPXPkd8DAjk57FZP2lyrl44+k
SguI68XJ+sScSS1ti2nhvwJq72te0iCYjCCD+fF4fKOCKy46Q3O455YmQGItLBOH
qj68B3HFQ4P7Pm/I973a+m9s+izFB/Od11MdZ6WGx97YfiuGENXTtopIYesr5h0Y
wPVJPHCfjzvtUc42baXrqrXngPYPHd5+LY8vPfya1vf18ZM3Ersqnjue69RuX9bm
dhKs7X+G1V9AMSf/dMRfthXxpEoL4xmo/JDEIFY8qy2TnDbFpQg2tOUs/K5dd+oQ
+YlClNp6c70ByfDy2EDVDnKrxWUMtKOt33g5P4wtgGF7fpR4T2TE+15InyULV0XF
lckS86F7E5yEKgaoKqcOD8EJrbmcMMtExFWaQ3zltl6UMI0sjeZ44YI/WJUy7z0F
6I/yVlpMrUStuUtdFNfK+1cWpnt/+Q+y9De5CWQeFJV3mNr5Z0d25vsjCKuvoOLt
BAY1D0kGNFihACmkiAF4EFt49I8/r8vBQOVczus5HTyuyt8GWHsMdxBUg/Nzakqr
NsszG1HSCr+h7QLbgxexXtNd7mc+YRHCvrHQJzn2d6ejRK570SVaaJVWpCt7PzBx
L+/+RCt54x+hMo94oQDyoxfnqiMnYeu9vGs6kkbc3tvLF/C8hzcoboBTCfsvIUiQ
x3mN5mTq8nwA0vscl8bjnGFpDM2iZVWWL67nc70h6REjur/yB1egUZX1hK4elY/n
sMOdCQSV+phiLW9h4qCEiekWe+vypnw4uYv0HZKvjqVb08MIL/PtRl3vphIM70p4
bQSqSzH8C6XqJ3KpVUQfdJ1Hs+fMQLeN3IoVMF15ZoArnRDNSmKeItcbzZJTiu8W
Mnhk5wL04J9yYOT49GHtUDiR43oFGpIfNQDXoNCQDokFN/UpiQ7CmZ1pokhKBcBx
QJ3ObkqbLfX3PcjxexTOPpwZc3ALCGrYX7u/MtF1MrbP4IB5lOhJQDFk4dEiTRCn
UPR+/tfNoK86ZfNLhg4PAlQsd/neqhxsnm1dQP+tmzzjXUn0580ivFCT8G60Hq8p
pvz6GQbkd2YkMagQ82EaYNODWPYYXikbjBrWg1Oeaowy8YNa2HZxwu+C90AgqfFC
qnZ+8KvpYWMi5lT8mlE/vuufx85ttQQcIxR1+e1OlXYo9YHxT1vYSJPjoocMm2tr
mElPMxQrZUVku/ZHn2zgHAGe5wk5fRBWWqqTBXFyIgenH7eWd7QXplA2iSUIVmgL
3AHItQtPPeT7gJUIeoZRfquDOr8WQjx4SX4sBdMlE5owTYYtk7vGY8b6q31hlk+P
OQniRr1dePiQGC6+W+PnpWEV7dxjl9+41iW5Kx74nVZdzMRdBv1Ot7LDXJsUHI3G
n9x2GuI9NACNRiWW8Mba4TCipvGkCUWO7iFsQ/kUplMMQWlGExs3fDUmgq/7WJoP
4yVdo+2EyAbgyp8j70rDnVEf0jcM+fw+X2//abM1hTpDFtu3AToR8oBHzd8bISbp
dGr8l8T3yCezQ1MJ9LbzYnDthnG0Hrfd/nfzUPbS+NUSQym5uRy9UYJLcFoU/0ne
LTOvclf3USjx2Zk/PfJCMekjxx9JSk9iBp9hpgwhsWx9MQJbmLcv5sOuKf8Qb/Lj
oY6q2ofZSM6wdEPDUcMgadReIhNpYT8YPZ5S6BFyTxtxMYZ8OHHLDTQMiKcv/rHp
gWjdiL2fmhiIBKRGMH2akRIYE70WOS6bipHiNn5n3xTs+/6e+IaVh8TgyLUfhK5h
Q1U6LjRGkjRRkZryjzMkgozjUyivd+uYTv/o7XyTXuFfIm32bUGaLRSDOaWB7kuL
NOoafit1Qqihy7AdMhx9BY2lf1SG5z5lUuDr/DfrxQdU7keC9QYcdrogiLbExeRY
/YbTw/TQncLg6Wyobyo+uBJsnIbysfoO6lVRc/f+oc8ApT+MWeRJ2ond5r/l5vdE
b0fl1CSrlUeg0qoSzimHia2hcFJhX/D5dwH5ocZ9nlcs7EeVWjKpsb2GIMRr82r3
1mEoE9MsVD0Jqatx2mffCV/Cja62wmHK8TOV8JuAhEi+DLV7jridi4017GfHtJqg
IRp0fgBUug1j/X7nsatXBL7iYpGf3VXyBJIyhgib87RQuT3o9SR9iHav+XI05vcW
0T7Hhl/Li8H9iHqHt1liCtJKQY5dO9XjnWc2H/dgwgtlKwQ7+PeDeWYWP1KcxjYe
yp9GQy3UBcGVQkgWS1+XuczoNLXuEgQybaJGvNutGBgKpCDZMGNOmiDrYESTzB+1
DYpbWDf7/e+3b99dfDgYyoZdfdVy+sAxrWryJv8xGlaanzb71XHbQOpTj2HbYnE7
9rwq54viuhNtp+eI8d+/eVYhGKPOo6JOQdX1sOzFNWn0n3JU7dOjCu8DR//bMo8Q
hrY/yJ0+a3wHJun59eDXQ2Bs1YB2SraZqSYMt/Iyt4C8lYyVbAU8u4OE3Q4W0sgw
QwbkRkNs4KsdmpgdYhki6j+jFM5JjWusyPs4RKrT5ZXZipxSiPWj5BUqC8iL8fD0
XcvMsVObRB0wkRYRdtF0n/19mBH0JyBlgDDjIGIMf46EuxcNEqklwPO43t9Sd9Yt
ebXoEz6jVdkaeT4W3WVvUlPDRHatAT8rPMkLsIFsBEHxBTrmAUraRF7NZXqirJGy
oGsHPEt1c//A4h96Vr/l35lLwoudHz/uRFyNJSHYF4lQHehQQuMAxZKI5ux3kLvI
TUVFONj8GHzs10V1ojts6Nd+VjaBP5pSCaKReePaYrNIEqwrv16+QR4eUx20Tg34
j0qp1iNaPe8r4/xmu9YF4vG9g2Ni8EIl5ajekgBXl5QworDSMiasFpj3UVWG8BFT
gidQyNmLQvZTT/MnbdsmYWLZK7X7Fpw2nL1iXx+G/mWPoHBR0oI2zzseZOqut5R5
MNTNA0aVGhgszMnWotMrT7eBZAbljDPhPvWbNjTER/HRLE1xcmxqY/8KjJ+5SCZD
wUUR9krvHcaSIONvWw8K54Zy8l96h6PSnfOqCG5lO7i796zsUKQxT5ZSLzzcNEB0
rKCRGNAMEfdkwW3riVk9e9QI9xIM3sONRr5JeoADGviyi1mlBJ/T+BuM1WH5tnW+
highFBhXQXsJ9QtRfo8GUnd3Sz9rTwdLISdm8xdYjsHudVRZJMW6pAYdgUwwwVg7
TjQ4BW5clcZJQ9Gks/90/C+H+7cdVYUb/YNYnexj3dhZIcOCOxqU+woTHhN5Kqa2
m8oyGFf8mFwwCfAi4/Dya9FOJeb3KPN8SEXdn4MRQLkb0hHld/ToGkljlRLPG375
HI3QDurjcdR1WZCpHAWf/RVTuB+PsUWETHYQseWWhOxEjWtYIaTFRKe2nBgCPjRU
jJBk5sNeh3TNY3kZdvqxI0zzqPe8F29/yhoyuxpznX+n4IX4tV57sOmFSuvqLPm9
tYThAvGh+v/Vlt/G55BSfJxrjGwjjYZe1MCz2lkYma7RKi8O1def55jZzHkI67gZ
NDkRjpVY60pIoRDS2z+B1UpBlp+uN/qEGWJwfbnP/kzFr40RkRrPbX2Gl2ShaWtV
jR0gAoEHxCg26qsdFvBwmdK0woqUColr7gtiyrbWQnm01fclgTltFzfrfu9rwdLV
09VygndofXTeY8Dgrw7HMv6ir94b4W0MLHB17kq79e69FcA1eavTrX+qZ4k050tw
x95gfEOqcbupV16Bbp4FcZwJ3viZbiTlsUUKW9WdSszd/cq4VZ+uxa9HwTySsVYh
WeQR49qlxXMmqG7osdpjpsj0ep52qpcMBXhMTRifk0tkXt2r/8bDIvkm/5Ozkx8w
YT3i4PjGUINtM7ylEVELIsGde3ocfbvSae1Y1naePn2F+LC8j8BygdclAUTv0yoR
QIgWj4IqRczGw2JuixdjVP0BnfLCeax5Po55WVMDIy2j0q4hLOgz8EyqkpOx1y6W
jBF+m1TcR6FEVFPc6BI7VWctoqeAX6tbq72JJWOf0IkMT3EX9+XiX7gyh2iG1fec
QrSvoUKNPw55kuA85sOCyouVZui/uvEZOZyQpn4jNqn8wQQ0ByrApU0jnDEbwknm
Uqfj9Wnm2GCOc6MngVPc4/Qt9Ov6+QkXtsgKdfGM4Cyq3Et7xC+4oAlgvgVSO62y
QCvs3kUjitBYaN7hyFWtMDz36mwQHvzRZSwEghXR+F03HRNQ6aVSmO/D2DEBjUG8
mtC7X6MYdG2NO0VuNhGRStJW3CstFHIylWdyu3KqwX+iRXeDuBPkaFRY/6yRWpxz
SFA+xc+5MIPhDKUu3wDf4b2cGXRhKZ5BUe376UG9fox66gxWY6uuf7C5gyGdM7Si
SwumQp+cIRQK+bJAMYLyqdYkeTlwvmtiSQfMSZ6KgAg6PWCQHAs7wUVY7Ec8RSPf
YrWiAi7lHYkExjncvivfV6S4x/HbIENVt20xrGNh4bwLVwWdWFmSArBHjnLXqCI5
LmUSI6fSyGSBhWb6c/zkKuAwHj9ZbSejXt0BWYT5ryxlw8zgkGGvoSx0BccBZJE8
wgTbT4BD2jexvHViKlqTOUf0SMVnQ0nhNoUF4HEAIoybQcspOEV/8feMmpOTT9Et
DwbaZbU2V5B2ECfhjIFOuAaKc+51bDAYQCOH8boNpYPB2+Fp7DAlEeq9bIRKWXNY
i1B733tjD/NixLetzZ1ihwvN6uC4LdVIwO7XM+05GM7eDa4DkgqI0JoKFiWEgzA8
deoPEsEedpHj7elX4APBUgxAQ5ahHuyOwhSnx18J8fcDizIkE9wk+OHliLxDSYuv
xjYKB7k/NFTxszo+SZ6vwY8aFEZFmZD96mo+MZfvBuv7uPSLFoFwNr4WT594QZ3t
2A11F2R98sKhrkhxWn7Q+C5ub9vaQyNPA+XkhNVLlX3WxHrygRE29i9cXaKqcfcc
v2yEPH4VkV4Lv283gV9KeKloPoDGCFwLCKh78oyGryiX6k0SIFtvADf+UOZieFcS
+8WdKiEAzyluuaIjrVbIRtRHQ3urdknRL73i8HdYZfuX3RWoOTaROf9kv27N4I4c
jqml7nnD81LEYgFQ18zvl4olkBjqyadYBeZe434dOdBA2fS+uZevtlsplIkYpdCb
zjrvwoc0ihcDyeUp2Rau1J6CoxPfp/N5BZYaEfN6DRVvcrH5r0QuNjerPMERQQXp
EX4CJLx7aDGm3WAbQDYGZwm5JsoI9Ad787ElRP7Tvy0+9nr2HbWBHC5v8GDUW8vU
20ksesDpMAHxW/VkZ0caDosDONFM36PTqNWEp00Yaug16Fr+hAQLK8v0guSWCDsu
Mk7+UodGN33Aoqu/JNbvYfLWttcvsYe5dZimXJzQ80ulqP8Fu8Q5vbFYHyALoIRi
OWLOrlzDJzR0+izJ7POPrpxoFx896c8jZlwOL10ZxeARYbRZQbAg2VhMWVNC+Z46
SF/lZj6HymX2Nz+7dFY4jsLzsDlXMF7U+vBzNcnmILzxevyDTCV/hHq1EMpzdtSM
XFgOxEnbhM2x/lyGJFoVzxqV6a9RsCmRWE2Gx1AzIcI/dJmqDb6AG23gpOhYZPtp
/jm4BzPRExh56VsVfzYmCoW+THI1UaHjTR7VLIjYJikhnAyUaGgrj9fEHmHsH/xQ
5t9oFg5J6Ma2fBeYlNb8+aGrTopnqZJ1DNgkc6rYABdNK8RAfEqHGX/gIyLKxA3/
OfmgFhWDMlyi77QSsWr9wUgcrexESO845hLsJ5Fyd+l06w1wUNnfE4Ypy+YWmhyM
WPIefj6CLLPvp+sjLbCOI/IWtIJu5OSf5x7NxS379tI7cdVrItdzt2Nh6ysxYwNr
otMAMWZ0eyvni2gF8vbTFc9hw6YVh8oMPj0E/oE9bpIpmrMu7/U6fio5+AcDkFoz
A6SnFYXo1iAMYMKdDZ6V1j89/ZtbS+oupn2DV/bfzpNeHmC2WZizjx4aoKOnTJlB
xiGPcrrfWRaGEFoIuVLtO0VyV4BCKce7SaLitYziztyPJqd4EYjvcafbras4zO21
X8f+rr1314ZN0agxX58ar8bvBfMBxdEhbiO6mS65ju4uT/r/BgXiJ7GqRi6aizJ3
E64fV9eTuosLcU5ipURjgAJCOc2DHwC+bGTZ/+QQ0VQDxdCBW5RMc+nCUIYrI6rT
kmEMVseNhKtb4zMqU87NVVCMVIsSSCftxQlZLcYIIf5u34z8aiE0SHAHXit1CzjM
smjOvV9x9mSMM+7QlDekuRznX5ordJuuM/0NxLyytR8r9oh6u003inhSrJepaAOc
n1mfDOgKjXqdW8sHHzAKqNfQeqbwpJdz9m9Wc6LUGcJUd3UnvlPnBeuFc00iGKaK
soaT71rU0d3Ahp+8SDw3PIX1oemX2Tlwg/wyFN0I1uRd1eEqrwVr1YuGtWA7DZgG
XoHRBrr8t5rPEIL/FdJa/E5ByNwFQiTDUv7EOx/CqSfrXd6jAf4PXT4GfeJPYv1h
o0JUXGlRZ/0C7uo0GttYLI91yIGHd8aWbBxAvEHbRxmbfFY7xt3R/eZq3+BwFe1d
SlzWTrXtAYCfyid0+jaThRXV2sFm5FaKI3R6f5+oQQiane7fGiQWb6AsJKLirOtN
qbA1oKNAYIlTm6AQML+ff3FvE51ReSx9u1h10vCFyG9p+H/FSm0Enc+bvmtgU02o
JQanG62micoHnb+Dj95m/a8h1Qg/rSVXChxFerA32UQpJeXYrktZJRlkVTF4oKZh
NE+2+q3XomhhZZRrEkcO8sKE22pZus+VlP9xRZwwkWvyg80roG6Le/6Uvqf5CL2v
XcDbhi9hFu4oynxQd70LtIyJ6oTt/UQg5F78ZAGk3XvDUGJgN3W9iuxsfQ/MO3Mx
AcK/+ZzUmQ9BgUFA7mj1dGTjnPJ+xNm46BSW2O6aqDcXUcukhQ+JXOWfilbs9JCG
ZDHbJH70JF4asY0BktdeLD5GT+m9+zmYIglY+T3Lt9UHBIKrwHcpTyl7MynGUCMz
PmyBEEdV3NsqUm60kzemt6rw2t0vVqA3awRzqRNxWr8uq8qbSwilYbFg14k4cfba
JKiRvGYNchO89b5FlrLuEExcFkhNYNBjsLMmWPpnQkpgYvz4gDS7lECJYQrV51sw
s4n7FoE0XNh9S7PhiEp1eDdFSXxStyeJArwUicAfIM50ZolvT5dHhs7YLrRs9Z4m
tGTlbCH1gX7NZl6Yx3R0IFloRdSqdaB36SZc/Jtm4IbRFjLNzg7a/f9E7YVxFXep
8Xpu1/QBn+185gPZsxWZ7qe3V5vVQvVarEEGc2hjmVbbEE56l5GbL53YNG6zfCjT
PTG+LptVRKFyj5wld/HRYEr4ht2OWrwh9dzXH+0WzYAjrV+alt1ah8Gmus/GZ39t
+pdCZ4kMMIxfu58XoMQYzqxMglfgTFP0Ua4b0eNCJf0Y1WbNPtADyeyleO0FF6DX
k2Nb6PLFuyPDKcf8kjMbs1nePKSFuDfLbYWObZoo+n8uKC31uLTjSZgZvp+DikDt
NFAtFtGOLryKi5//Z848wbjQZqkY0B6PMZ/inOX+NMPC6uAf5NPvSe70C5ZRujP7
7qMFLe4c7peO6JxytlA+UlVy6isFEkFudBZF3lU7cXRJbm5CCDESTY5HGgubBksa
zfKbaMXL5NSLEyJV2adyIsw00C4TS2CaDzruZsKqnSjpjNJF4OaIb1xjZx6P8I/t
H/lZ9TJxGE54LXzTQGOCiWhsSlp5eix6DWMYOc7wSNRxBfdm5C8QBMf7+k8gH7Fo
SBWwoyaypPLJIFkx0PMEUe7YAkzG7SSB+MPa+LzzBP6PqNOhhA4RvGXCdSi98s9D
zkAYUyIa890q++9ahSorllQ9Rd4jDscX6ctGHEthqmjzp10I5NYz6omkq9b/FqQc
DggiLvViiA7uZMTEe0nCgoOGfoHcDjpo03RfeTVGkWWuarhw6dxPRP4t+D4eKqPM
3u9HoR4oklqOKElqQ5PitE/9oD9MlbQEPhCp26IkUpZvVYL7vdFBEI8YSyux7K2w
xu5i/+W8n5jnldF2oNn5mX4tj7hsRqUrLPYj83VfBXUSCn18us+ugf3quvanR2my
3ggKjNGzPADgCP4UHqzg6BUAcUMH1vMBZJ2MMDGoVoZqOWRScNd5wtdXiIhgh5VX
YDJa3kr/OmFrXOA6lqI5D3NFzE+oZs92V0L4NsJMFOo3GjVW0+5EH+T6auf4OWRU
98DGzohMSl2UB3QZPCMO4gTDZzLRLuBAniynqVNq8NrOTdPNOXN9XVYDFJgfakLU
LjM4miRIBl1mMcTaUIvLU4ODAzMcBwefrLq9l85py1R/X7z8kDS317hHLgiaIJFl
bZ/5W8srXxrcXdCzDXnPcC3KlkSaOWjtT/1Fm0Nv+BKf3fLoqMEoUgonVc/Y3TCN
emShERpgjy361QcfEGnAgTbP5BIXbHwH5+LaWTv75huYuv1/2Ruj80YPiy5bngdH
PGjKjmHe/JXWuii+uxAofI74WLWiX0MVqOiT+YKloZnist9LmkasszTgKNSWJlwX
Ai5mKcQBJ8j0R0Y4snO06EPHbTNP88eerfz46dAWtOIH2GGsG7wrLJzYHTQrxbSI
/6fO/EihdtwDm+dxleH1jzEmbzVwRoIiqL15vWEZEztJp1CnWue2IsurYB4Jqudc
dR2kMDqnIewWZs/VqWP6kDvE/D4957BtOYew6OiDogc2gePC5OQZyImvWZhy2Ua8
R4/i7s7/LmffDhDf0jnMTjvdQORdhf0U7m32Nc+t+aAPrOgb2mDuFyDN1bqq7v+W
uilQVOXgG/9+jr1TnA8i6xqwusv0Us2cMdhshup3bVo4eCeDV8GEPntDieuhqqvO
wwgE7cAluD7E9Y4kwaMGLPmLUAuVJIdp/iZ73giUQSuTXo46r+P/c/aS/3zdvNGX
jFRVLYyiJDUWVUx1cVCLp7h2agn8bKtwxMZjgLo9J68LmErffoCCFM5JwGQG5Hg3
do1MGSu4BoQNjRK9IZoo2nTbRS3vjgTjps0yhwwjyTfvj6lLcchYEJB5mvgLgZhj
TCgTrf5U0jQYJjNC9e2fJQoG3Sw17B+NKeKh0aSo4r5IJx8LovgSdO6Yz85Me4Ud
OJ+5ugiAv4/6cPvM/KMRw0ixqs8Kj4iarVWRTnYJlCbG5c/elaA551q5NtAdcmms
yOi+zzjC4idpALxtbOIeebJsMWO5NqygF2A9/keqxNPMEoJP8dIhW3o4x8vWkODu
KMhxumZiKgaSIWco4QS7AIwQgA+JffaHvNgSvg5khQ48ES2cz5tzr5EkvURKO9Vx
3GilMDcMDzUij+2b3KGWDDhbeHZOc9WhyUUpeDt0okNBap9EjKcca1xa+1hLBdaO
ylk46jNh4JOW2ARZuA3RCvnKxnMBPtd4RsGy4SgByurdnsaedPE2nCqXNBP/bdrx
EQISIuKxg+frxWOlTdC9qUmmPHPDi4365ooPk7yumC7Qq0F+sW6yLha14jqU30zQ
fLgZCXO/YcpxknHzuLbi8wzlq/AzND9ffusBOHbXwfnPJZU7rCE4P2KkPxpy4McA
yrOWtVM/3PZIZVE1ydkrQhZrwCfOZmQT6Uw+sf68rZwe8kaKs5yqI4rr491BSw3o
/7tfJG3SHUu8ExRu1louAj2DG+AHaCpK4pgGMYjsagv50+kZHQ16toBsXVpGcuWj
5YdTRoBghJLVuNG0br7jx8iDeY2XD7o0mcRsKkqNAJCfPyVUKSTaOuJsNIqTxBp+
63iGMUZ94AfVsJ4RCa/pZy1uniQpbNCUv/U4Gl/u5uGgr/QlzieRSz1322ocx0Zx
97rMcc2VdSyrIo5zSqdJXd9qm+e6NAJ+AG+A5x1Y+q0oxZCdOWjO7qxRshGjL0iL
Wf2lfbqS7u5WUjLpgT+yKN/tD3f1XyYX+13BF9FicjvA4cYMRaJyPIMkuuWx6kcA
PeyolTi9bI1WK+t79d2oQ099hwJL+2pngRLvb4oxxACUF2B7xyW0bJhGxX8W/RZv
AWe1YwAN1cSJZEO5BX9tZFYWnohSuNHm5csfQMOMuhtW9jZ7iFJ1ppP06+opGK89
UfXAVdu4ap8SFYwGgbhVpvfywBUludZ1tvstJde6AWoUFnvZwti0HeSEpSXfj4rI
v1tFVnjgY5ngC3U9XAsU3zmIMIojm2FkQRW7mziM+o97U8RAP7hJ5/V1CcXEZPeS
cNC4eTylVq9LvI4rY8vW6RqLSNz3mm7FfGtsymjUoSlWSRK2U9qMjnArdYgNiY5i
sjAWKTjGrbXJbXGKFTfNudvlKnLW+FgfQbsufYzNRZplOF+/Wo1xIStteDydasrC
QTfQLn5iEuxgeKL+EIJK0BL+OgaolqobouvMPPuELINIfDuL9A3D6/MOe3+Pehg6
4/j/MDRAiQOs37KiuB4IYplkT2sdDSMisjShBCBmxygy2DNRvHYyJ5iugOTsoNvf
QzjrgZ1o9t+5P/C+flQp5przyYjUNrEbTdev/GfZSrz3sopKqnXWmK24HJcUxCo4
aj51Js3RyAUFfXzT20snQVwSly8M/BU7jyj4eYQFGseAfwpl4RBSCcDodUX3tD0q
MiZs0d3JaA6OzU/In35K322ZNAzzFSkeRjF8kk3VBO/HMXPCxnNuDP+tm24u5tfT
5kqy3PXmTyXIVGlnoYo2T0jTvi9hhe1YpKyESW3XQSw3nzss4+Lh2IBT9VmqyUq5
vRKQyk/IUd1TEdDfRGWQI3JUtceSVtTetIjYTSTjjQQfjmDGgLpXcN2vYMYC+bYJ
W9WIDqN64P7D5cn8w5m1Z4w4/nxCBt5TbLdhS67uDGusacm7x3s+svXkmPagiK6E
mV3/heFctkEgI78u+EHBy7LL8AqSYUSjLqj2IN2ljRyjcs6oWaI8TQikXcFyD17b
sbhQHP+VURyq6ACHksuKxWrLhRHbT1cj6V/Pi+UGoX6bEcucV44ATF+cNmTnuBZZ
IFHfLVC51/7d7t6xewz5g1EciMi6JbQd4/07S+TP1L6XpMs4wVkELII8N/CAPg5R
nkWr6k8LFckptTqHHt670GoI+ja/8hpbNpI4TFwosfcl1/H8InSR/dgRKCTAkEfv
vInxB44RC/cUzwXy+sqvsiLHR0yRv/HcS1otJUw93e18L7JE75R8CBzXfp+D9G2x
grMpZSVNvFsr7RZxPwxq+t+9uPw1HY9fI3QNecol5mpwqMnRSSmwmo3GBaX2NL2e
TcPI4r4MsKx7BZa8sB58pKeMhpQpToY4GgKApzLsdvm9S+s366i0A36CxnCFPzwZ
G7UYRA1ZVYDRa7ZyqavJeP1KLhBsPqt3xCoU4YwvZBI5tkQ+gqNNQwV7KCGuWOPu
8LFApDCN2Y7h05KIzlJx1ME3I4Dxt3ytmnFchua0CzJy4fW51htS0KrtiDJjBWjE
uc31cyDKLjMNEXxpzh9jDXM4Hi3lrw1Jh7eAygz8n5Ft6cS4ni1qQ1/0ZXV6v6BY
nPCmgmEDkp32WPCqM9hjCfd5o5TiotcjL5lJ9XTexSm0LCcc08m5J4JJNGPjDmV4
qbKd6W5Nmll7cOpLMuHDjl6av+SMvZlp3jWBbozQPenl9fDxC8OrAKwdesxLay7u
O+GaTC3j+2yuhS5HQ3O8A4ZExn7Q5Ryrom5fjds9zaTrtW7bi4T5jpJfRkQsC2xt
3BjbknDqvbvQSkGYtUi7oJ0xR+v90rrNVFP7Whg2dqhPARIoRPeYCy9W51yNNWZD
GJv5dodvlHQ0ohFWd3SOxktWo8GZHaCA826crrQmaG75g/HXGXGxCmAXBv+/pk0n
GvhC+XoyFpldqeu39A0btyf3dtED988un7Lvizoc5HeCh6gCw7h+xOLFPG4nEVN1
pPG5yvDRD3Z38vQwTo9x7VoIOL5ec1QuC+l1JxkICX95odzfkFSvA08c9re3ExBt
iXALIndoew7W4BE9Y4/pMIKoEFpj9OqCkOXDgTqaV2GNPi+NyBQ/HpcRQRBCtdiZ
FYey1w+NmP2NG/5KvbEskpj/1ZSeeNi/ZPiMbLR9eyqtrBJ4RWj3BtTTBp0uHxYE
fpIXDvt4I1QS/a65L/NAsMneVp2FSPdRtxmK6smMMtnJoGTiMzSVNgACn1Igu7lI
IbEofjTwD+0E6NHHdOIZIRicLQrPe74ibqIjAksdH6fo4jw+A/YTTrg4cC0b//Ax
v7sgNSdrIMU0RftvEP5Ceox+YI2PJpm8SAd+oAqV4kmAla2c8GzVMpQATsaaMpZB
6P7v6jltbI6q86nUP0DkkgMperRNoVYqvQOy8ojpbF2VXdiEAWAzMW/hJXflrNKm
G6YnymblRdX1AoPg+uNw7tzZM3BLrnWocOkLN2gV/R45AgepfNzJfa0RlOZMuFrc
7FwNxEmm/7RsL7nnrBhfD1948g/2PjmOx7rElVl7IUaWn1YRvv97trxxF+Mva2ru
1YnLQ2MKZzhD+RxNmVg1O/MK9oPaxhkRmg5kbRW5sAW73h3J+lWxfNIxu7MLEJ+L
YmFxncnRe8x/NJJx7k87WEWZpvmLL7Ytx5vtSrf0QLYhuNEIJ2Fk2pt4sn50+dFj
hG3r9EttCu4nBIafEb7+E2wc2AaU4EEaNhKT+Xi63ngoXJ+W01uqFixh8B7q7bQi
gKYcGWWyeirs/JTzGIN2fipywRIRR/4CxzmCTMz0Pjb+gBDGckoZwtmHgeTJWyB/
hZjZLL+in7DduD17vCbco+cfuauqsKdR2LDBVqG7IAmXsn3LhEJ0C3Uijc6GoLxz
Nh1OHTe1rEhnaEHvPQIiuWa3QaTfjRocSrqvsu4jAIPBYoFKLMoTFbJzKaHjPkLw
gPSQN4ssWdjJshm0jqHCQpcufxbuhOWJup4q2jvE+7Q+/kcZXK8XjMfkFmSGWrTU
A3cEtatBXWUPmIlM7d+fMcX6YedOW+Z0SVLX3IIg3kCpWLOghiKF8VP5JS35Vh2R
HOLQkI1ufaWpHFGNdt2aF5RCiHIYVv8yQrp0xSO8i3tD48tzbIFD0VvaYzut3+H4
JUQAkYrzv63wjac4H1nEX/Ve3PlX1gEufV3UL1sX1aYQofyjyYzKvK+7JV6v+V/F
K+OjsTuvhATTOHw2Qc8vmaQo9wGij4uifgay9x4173axhNF3EX7SWQbLktuT4hXL
TyUMAeRlueG1pGNfYED1uXme0azoIJ1pothRIkWHN4k+so2BG/hE4RlZl2DS8zLI
lWvNCSevSiwq2YOsa8mjJgHxaC7dlVEI+Nvy+wybGQPiVF+sN+C+ClVGUrdaVC4W
enFupGNyWdLSkvh/QehS6eQ5itvS7WO3xoc4ip1PgIIRdZMyytfmXGRKEiv/07PB
fWzt9VvjK/BuWgWBpP/4+90YRnAMKnJUOEM0Uepf0Hx3iEHs1znJ5mpQ6hfDmDuh
+9ALNiJz9js+bG+IfZD5WdjG2Bhfm6tpcSgL9JWXhSm+k5DdfmbG+CxWI3STUma1
iZQsttlNh8IfkdJlv9wLHBVwfijQGew9XDG4fECJx8PvEILzivFgtoOz5SyGoUsh
EgIkPCnj3xUPD/8oYmMb4SV6+qCVdemlEhmCUg7mfrQVa0WJGOsE/ZeN1PCHlEnr
DT3eal+B7H7K+uU8Q9s78L7O2EvQNrWvYvwSGo91wRz+WToQywdQ6arDdy+pCgyY
gXhi5iXWzmd3Q62pqvwMq0WN6cnPegFxbt1bg7FNrCnl7vT3W1JvTeWvlr5DqbV4
U1i1yswjEqYbcXCJdD9A1aLjwkDG7NvSjHP+KNlZggzW17C3BjG7g5sPVpg7z1ZQ
ANouryagTGcDCaN8ebpHKMhZIzwl6aCDVvSjPipfnETdzAeiMv5I+k1k6NLqr5LD
3BPj49tdRPzQLFNfJWCms1tQ9zIqpTRY9vXjeeILopqUOqrpz8zxBcDHBRFFvdaU
MOvyBay1kCLlTOZhS+gKu0rVVsXJ30W+ST09vddc/Lqx73fOFn7KJzNHCEe5XcZz
N1b1WjKFC4TXov8v438pkm85GrT1258WJTvo8r8oNx4vUeW0Bhc2AUXQNQZAKouL
/X346gnv5iOKKVXsm9f6KQBE+IwbJup8nl2PpaqNv1mKQQh0rYD+3OiD73PZXlXM
vNa0hBjT1b0fCT0yzhlPfnwhAY618QJaFxwYWcM1LvLqDKgW1DI9aIaEQXQWCBDv
s5RKoEsFTZ3P41Yym8Aiav20/vU4M1COp2vWMf1viFV+3FwjK72IOFtMz426qx1w
B/TlA9HUvDUTnJKlJl38sfMNaI1UQRdbQfny3VaaO2UFLPYm0CTL6UGh4wbL2R8m
idOkvQO4pcxdDgVMiiMGwLwIYbP3aBS4+QbJv8VIVacUKQbKaPi9j9o6bUGrSzlH
tRrUUECHGUAHEXTSeIXQjrRsmoee79ATIWNMSdvJioLoneQ/D+y9A9e0Qwe2LsEP
wEDaR3Z+vTuuqGa/tyNJExnWAZPQJJc64M6zVWV3IL5CgnwWNAG5NT6hS2o2N22B
MjqMY9gKAmqA75NOUGDrxVBIPxeMsz4EGW7Oo5q7WNgmV3xTocIvj0/IkbMn/Qot
me3NG9ZTsdNpQj+YIKmZ2M5TIzc8cDj+AhYN0MMTaGUOHAfEo7KQUFEVg3uZXVBr
OgcCCEaOsgy+wy/giDNAFn1PE0td52IQ0hU6nCZ320Y8fTdyJXTSU1mNhKZC7E6o
cW0H7YJNBW1vDi/WvAuc1hK9wVjpVRWHDS8dbqS3GGs7xsgHqbYmo9Fuxyp05sYV
I/5sRiFRO1i8k27A/4FUUj1TiTL7Esa/dlcpw26JsmQGpLf9BIC6Dl2hGKCUnuPl
H+ueiQImwroDDsEWg1Z/fkcnVt1toP3jrt2YzQ/zsSibNLfwl0fgjO7PThcIcCbT
jfaUwU+PfuzOVinBr/bGL9m2P1Zg+XxyDDdoivDxeaKTs5VO0Eojmp1Ps3HncM55
c1sa9SynhgSNw3HyOxXRlAMOxuITrEtMS0frFh3a0URdPkhw/GQDuSqFDumHtJoS
qETX6jiSVpBbc2hJuCEjgFK/MzFA2H5mt/B8skYf2vG5XG/aVb8FGGWcyzrHczbl
bLFozwCPfoRzCOhMVfoVd592QPDp22W+//dlUuWG7Ttiz5SrGFs2Sx+ibXCZx+Kt
FA6AZR00nBmErlzPV+Dr12eLJAzqyYSO+1HKtb1lk0VfF8yP8TEg6yuCA12KzZJM
U/lv/Txp+GoOcEl9sk1wuUZRakzKvQUtE8f3R4Iko76Wl6YipnFzjtDLHENGSK5/
eHJXvrdcnxgL++yfp4m6sGEebrbpCvp14AWf56IzBiMkStwl3ON0LAXTTJ/ieWAC
P7dgrThkhhgoYEp1YyHsKN8SAPqO2ZBTT/t3pG39GJyHbz+/WEa3PoJp26jZM6by
CA6o1WASesFmBYAwAE/jiTuWywRV9bU6wfjknek+76vHaQc7jLfvtcglW8Gg7vCk
e8IjzQalgi2+FSRDBbl60nYUbi+Igg7uCuWDTkcCWDxk7lcAHvODPNCGUXZRPjCX
GOExmEiR6l+jl7dKvGgvDrTOihv+khteHEjwifFYwL/+td9xqE4FYuDtzqxpk1J9
QKEUUbqz0ACBy4Dcn0fD+0TV+lp3fPOCc5dpU4m0aGxH9ge8hM6++2jUrGYfb7sT
b4fhWT9xFEGt8nHs8GPZ2Vl8WITstVZ/J1CUwtQ7juTmOWafxrGjuqDraGA/6fk7
MwbfVzYIDL55SmBRTMtG7uqm5N28Y0wrjqkfkl0wJ8IeYxKDO6WVAVSjw5a9cSWa
b4Qc9W/tGrjzCLsEyBvAK3UcSGxhuqBh4EgKFvVDH+BP/5/g9TY4zu5RPUvH4aW6
r/olTNX/nKwK8mWTff976sFjP+U6aMnCQGU1ty28RDic2wjdVLW8i4/n6rdFGrb8
9uHq7JSVLfWYt38N3Ov4vQ0+fd3zr4T6LUe810NS6s8FfzlHJkv7/37X8ra2gCsx
8ekIJcMn1XXmUBwWzLLfIufC2JoEFvAbBg2OBkrqVIcyWePF0bFGbKo0jCroky6M
5eTdVhJPGSI+FcZMljQSclxi9gmKnd86i9U5rSkQobD1fN9Yns5QVYkomzh+3zyg
RCj7GlHy5XlK7RYJHGBTTNWMECzM1XBxGtqlW804YdUb+Fb0v7jcHHM88Mkb5Qmm
lxcc4FWhz/MLHqPyaoBMzWp+ca1xcXTEN6EikcpvWe1fWYHe+KYjJ9g4NTJGPfI7
ccr78ieUaG0oBTGmns5yADtg0/UND2NzvhQmoAnUe7BCLGJvX2rQ8P7ljYi0M8EE
SDfwAqZ/7qM2HtWmR+jau2TLbfNIyQTx/5QP/T3JUVsvH4C3xLVwT/xqLu618eZc
qPv8O83LoOUDJAXocrofp3Amcc6IQlZ+dM7Uh0yfZYpU3C9+HxBt+k3d/hmKnmg3
iBg5xt7NB9YWYbj46wroGAaKmpQcFJ4epAgYwmSWd5cgQOjLzwzYC0hFOBmpQUe/
kH5mCIuDs+O8xbvfBWpfZVvshSul4pFFDDdTi/hjOt96h2UrucvpljywsEtoucot
OKXVqRDZ6jgRcvFJHjM1hQEAhl9nbFHeMuM9Hf6/d1gxdjY4s/MObT2nTBJPPDsZ
rl6npD4jNM3Yf1Yngbin91ZBnO3fgL9zvy0vLq2wo/9fHkKJu/TVdN28YtGiIjJF
nPYKohwqHF/nT6VZq6xTDTqhExculW+q9VzqNlgInti7lZwq0Tn7fwuU+9ZrwpTa
LPRswkLB5svZnkbCuSTdtQe11QSNblg9njoKwreGmPKAcMTyjz2bY5mHD1zsHoTW
uyre1IdZNyBXaWyOvc+CF/wrZzDGf+YJ7nXN15fuj4EzCE083hhqyrwYWF2UwNKd
Mhvg5WIJWKJo8J/+VhZvOx8kx1/pvNuCGBKMgTqtMkknjjc4H2UZh9YQxsTdav+m
X2trDAOH9qJSZ9AYD/NVftVs5GW/kC51sHLscRWYr5IrJk56EYtWmWcE0yDU0T0m
x1eAdEOXe23Y3Nqm3wM0JUeavxVp2ogof+4iqh5zX9DA2nd75ruuFTOGji3nHLVI
or3U12IwyPlhdtpRO6/GmmrUhs0YvUCz4vrMX8MWLNmucw7E9OEusMztdL7wvcKT
s5vTK/DXBXStONniBUcK2c4tr6cGmNctbe9xak5ljgie6DHAUsWvNY3vn/J8Ofq+
jkjAdLHCX8HxV7uHqMeFugZoGHR08qNJjbObJp3xUhjeVDgAYy3EJ7pdXMXdigEv
KH95iv5oc2Xlb0MLXGtYyab1I9wUxyoy2EZTIuV0untPrkEmrR5hJOcaPbg4W1XY
x665WVdPhLym2owP7FjfWYocqBldwT+3c3A7upyACw+FQn6RcqUKm/X2Hlfgz/GG
C+7FHi3Ja0sMXj0D6ZjNwTVmwEZU1Ja4xpEP/ttdV6uLidUPUfIGL33jP5scPjqs
C7vSEe2otZvl2k9Rb7rhFr/ozVZ1yfVf9ri1J9s4IVqrDjtQ6gRBC/f6J4Ticloi
4EDAO1m1BTk5KGwVYuyjaDBHOM2pXplmEpYY5t2TU/DB1iBN+psPGAhTej4N0kfO
gSIrvWhrdhAlMr1dJiE626nHnnL8RjS0hKbsuah3bkudcP6IK12WmXAidZ0yco5s
/AP6S+o/4M0dCzicjV1A46vU6F6sQwIxM+WqfMRgRde2UrUpJVttApbNZvh5wgcW
kLRumtepKit0K8x1tzGEd8Zgw+7aKVrJTMktP+4MABVevxv2cmyvOqtvjztnfhQz
lGBMiG/GUHC07UfVoCbp6b0loG4h2s5+Ch3H3SJ0sv+XMTrTeEFvtKA8p3hsrpYB
EyaJGjpTuyD7Oh6QjypflQ1jW3+LlunlrmVVyjnHoaA0+DneHZyyC87gY1mvQ0rW
ct9NA25iwBSfOycZ8mv8htTxj9dH5N4xjkHXRpTtYCevSphqNrUyC2jIkeZMGHcE
WUMZGAiV52zMPCUq1sqezQJmiPmYBc2vdUaL5Dc0mgUEEYqJJM+5edhCNQYkZnAi
20w3R3We8ia5zhRIxSb7L+JdFCEmyTQ4YTLm1oSMlP/bawmiNjgJtwKmYK9R0Q4X
LVbds6sB0igaKRUDUCnqaLpcGKdDJNBNjjn58Pci1SS3UYw8bg5bFeJDxzjRV59L
qSHfPYtNCMzn3b6YqsD4bPFzkUSufxErH+07+saBm3/2vUy22a1lmbyYEEoz0sB5
2UtrAkp+kD9J68Tp2m97LlMQ5YC0LhvjTY/wF55l/ZdqTjUaAM4gCRW/YFosdek2
9QWVet16vCX+YWGUZKHDs1dKEfrobhSNFOCgUA7e7yWQyekQ6RlHmr6Wx2T3xobP
oaflUO2BSuAJTThxHG3h7rarlo7cpCdJfdi3OSZPncohv5q9CjpodDh7JStgPGWN
Zt1PCbOPsL8AKeVNjvuH0DoSELJTahEIXiDrFAhq5xKiYhNZknIvLRtUwHEIWOkH
LJJYgDa4CixnNFyoKmLSH/qzGS9ZUKyEvV1m9hK79tkwJLhNQkkua6ElcCc+O2LE
nDCWzsPLGJSIMIwlJacewzhrrP1stwqY7zmH4tYizVKJ2XBmYxLzeq5hjF0Q6tmj
krK1eu2DVxkY5fYVD4qIxgHjmQBZSOUmi44EiwmUlIoVXdL/q90rq4WOdsy5psEG
uqSAkXC9kLyjmCyVkDQWcJm1aYOOSrxk7M6Jk/2tUYmeo+PIv/4ZBJ838dH4XE7A
2Zz0cNsg9OM22WB8ZJ438vwQr0sw8++dOC3TxQzR1adWyrBPVLUMZFxVkhbFpZKg
oQjUtF4H3o885RH/6U0D07fYRu8d7Ci5Bk0zYj0OdmQjf0Kst9KhcyUEfIIEJDc2
h3a+CFcgG1R1R81my/sugtBgPKxA0PBVTKI0P/agQBeHK6aA3X4IByjRw3cMgvXn
ILzwI9Ks6Kb0DcCwbMeEhCagUHzcCYhgzVPFVnwrNQconq1IZT57qUu3OOlveQS6
TrXgttAG1qD6jR944LusYdyjMbns7Q7UHgLKO06bBbQZdggxxSh+38N11a9owxYk
n3TigNbgLSIg24bNjjeM0uIFmvDFSU9VAZR/V0WFwskTZV+atkhW2iH/20UHpzOe
xFfm9pBs6ypb64JKADvNOsICNVIEyouvXY8VlMiHdiznyDJzwfBA7jmwsKU0J8Dl
TS1KmLudu+VfMd2MZhYl73MrUyjbCvSNtIag5lgjOzpeUIDhYgbC7aZDWNTlMUVu
WXrVyVwtv9dn33lQTjz1XoetY4L46GaNQgyxASoYW9WbFVFR4cI4bHMIJ5Nbjidz
uD4ag7iGVK2NXDUskuWHL8FtSmCkx76nWafn8sMJP7p9abeko8ma4oQoCbWpeueA
xpYpx0XvZf6VLy7m8Nl4p0oNoSzBNoqnBJLRP5Ur/m5mvGpLRZdi6S0YytrJRoZ1
AFbk3eFW+tIDqRPDCSKXlaB1bJ3qZ28QiqnZOduhtPKmJ0GGw7oqR/pexGDOMYa+
0vSjPQnli8Af1vXdbtFEzesHBNuyM4+/MXjVzGRS2uQq48m935g4Gx/DUOpKmaQ1
CDjCCh6wwMSyXU7E8Gi7oLrguuykuSlHc4S2PvlFMtsKlNgjaazOl78TUA+r+ToS
aay7Ph1JfYCbg8Gq7exFP6zEcLktqgKd+3kDLa/dP/wLWvGQL10ThHQ+TBv2jGpP
iXCemAEBsFnTOPu/LpA/AVgzV6OEjTPmdbcDCp7LvLUdEAVw2GSqsBnXjN0KmrwE
TG+YFu8vXSanGTUAO5g0LzuDGtZv0HkAPeDgoiyJH/Qa5oTCoIjGVStMYverP+JE
S7BQsPAQHhmC6duDBZbgEfFPC3mDwlX+IS7s4BTqFaTlqaC8ZwUMg+b25UM69xyI
7gTRWlI5Z7/G5nSNpu95jVEkWrStvkIDQzGQ+Dw+MTA47gL0iFLkfxJ49PWfCQCS
lQkENki5JSiAd3KdtEX0r87Qwu3q5XDrS5Oa7nnc0KKhhQijrbenjOFuwBPd+oWy
pQjhaVtSBbQF/NaM2el6XUcyy3gNQBHNgIzPVzzAJ8k7p8CLYpyYZkF3SEZHfguu
lgWMxSGybnqld2q28lW8WdvmVDbvkUL78RRjPpXgh/yAOO/tzUgfNB5HrPgPLpUB
VawikmVvX72XgEn6adbG4sU/FGRp88FrJr3GGb9Xz4OJFS5bXOfPjafneLpnBmeN
1PaW2V2qUwaV+LqwbkkzWLZtphrAp4l+o+au5m1bUNva/6YwFQ5cKvxPW2rl9+y+
6O1GExCEoPtYFKQcpwFGmnbIEHUaWPJ8LfRVZ+KPTcivXA0i8oKEj7/ifXBS5mjR
3RInDGSla2rCUqcsNFiNeXudD9xXwJHa663mHjmIGizA24lNmCJy6HvMf+vo+0el
XbRpW3tFHq/sRDFHSe0fKi3eFBI5MyzHmX6J67748fmjDUVQo99ScirwLxbgk20d
+I3mVgLptzE06JE1A6BPiEITtjQNVWhqvOn0HWVbKKtlvtfDbTA7hTTIVGQhFUXu
0dRU6LWTD0+zrfgJkv6nNunmYKrsNf1XTMF8dZsLsicGleEmhfqfp3AUxCRKo2Nt
XqWDcZGbNGEkzQQKBizRfPKhgShHDa91qRCAIX2VIvJJ8hgSl/Js1ZUJvKal+ZEC
LT/01BXdROd7Br6Z8oDwyWhzhF+0AQO/kUe2d1xUdH45h0c1se+CJ6c/0FHrK4Qg
hP7LHTZ64vTNEp9lQ9QNJXeW1ISR8jAU0RofZdK3ULEEm6IgrW5LN6+6WRoDFWXV
/FVFya6uKwqnZ+qA3+QeZzbA6kLHh8BaK0RG9q04Lli/b7FAGp7WNgzV69e/3Wmd
R7LLvA01gn4t7XcmUoQ3PEIguDqmu57Bd2EPbO3IcBI4qzJKp7kdUkqfqgHrhl8Y
g6oAPf9GYVz7+eUg8+xY/NlfufoJdNq2h9jr6LINe4T/P9TWd2pswFpaur7hu4rS
LBh5v3+d6Plao3XZSUAR5lqO9mAOvXk6k+hqyNdZjNal7VzAwYAJEPY9rgRSlgz9
i/l3T8QVRfoKrSjlvBe/nlca13qMpCLMtC9WMDSd5ri4weT620NJOL6LBdqz3iBl
fUmt1aie26Zg08BgQIF6Tmr8bchkZDco6HXc0EJo/FKcKSylDHzRKObdCRCFMyEk
9nEh2WQzhrrLxEL7RTx28HyRoEvrv2k+n76AA4tBn7kua9U2v78QH+l2mb3RLhDp
gBdrjHcG5boanu1ZdCakdLrBSX/ik49rmCN7FY3PH2mntIUrUKgh8aJd/TbWq+U/
1+tyaxhDMG2Ft2UxJCG8jGKM3NhgHxuJsKjFz/997115K5tp0tnMm0fJLh03cklh
L8zSOqac8Y2n6XGN6leJyf0n37gK+a2BhClfl0s7DEa60FvuKaqIskFiwHb9Jomk
9FRfpumFuZDSrm12bqUiKgX5/rtbb0Nd8balbOopb8/EJ8W8ge8Y3cMapixn7Hx5
pmRPx5VeeYWnX4yXNX06ZFX6dnb2d+tOXH2eRK7SVL6/qTet8HObzfKHtbGeWaUf
CB+CzrKVIb+ZPweQKB/QMaSmho7cTH0AaEhBDJ1SX5S8PHNdc1FBz+or5gTPu3vA
LCh0MwgTprdZwfG8BotXm078vHRZYI00IHdXXrDJYosbVbDlokl57zgchIZDgkFf
T3pPQ2pQEh8xWt8xnjE10we3yl21g/Uk699/CrubsQWwakrPT+V7sSH/THvbBrJC
KIcALVJdf7ewTM0xOEv4pbFi4KrWypcQ8zHK+HbfdiUa8Aq5iuqSTmaX+7BQbhar
AxMhmypXTP1KRcqEcRmh2WhASYSCM8QA9+jYHOMf2GETVbwgNfR/1jGfhUwY/G5F
YDNeXRtpRRsDYO08TqkDrOFdMhcaBT3JnaJKpB0Dd7esaxHDxk77g7WyC2d1BGzy
PePd3HdIMLGpckPsh4ZfMGJHBeVJX+/Lud1ZhwQ0a9bNJbGE2iryWDBCBqx23NeI
EIqlQLXe5Q3rQudMtVG88NOKtOXuMdbo+oNFmqsRr5rtIkVPtpqqw6GVLI6SmA1i
gMg5MXH3quyscG1eVCrN76fjMJZXrGzW7rTqg1YUiUqcSrHxoDjRr/0i6QoGghZs
4UmzbvnbZLxQHXUZM+yUQJaNGZ7fdPmmgfkgLnruvSwLOQWYft8vTrOuBxaL3Kjm
L6M3KhvCdbxykjaCiSqjEYwkxybYx/vho+Mz4E8zlPLL+geRf01f3sQPm3Tacfol
9ya+5ik1TEuPfGUHvXtxsRkeJ88+aC5WodLWtOM9wneTYcikxNBIwh+INRx/ZjsA
/2O/Sm4VNAdwHAIUGL0+GGwcP+dhtye4rgwKTh6tXz9qnS5/3IsPyxoIeYz/76SS
zZTgN0icyIcTqcCbmQpalj2MWsuGYhpa+lKbWHd7itvHAq4tUmxrGT/zgCdKOSuE
Yek8KjGaRB97PG+jZDGqbupDNc9+9x28LZ0o3TztYa0vM+NRJjSvqv4CELFadbw0
31whtnrYG2fh63BUTweiheHFY3cFatrrRRWslsWgfccQF0DoSSnbyVkIeZEx0sij
vgiCtpBYT0O3dav0YWeZKDnQAiDbGOkdXAWFw8Wr6s0+JHzlOJNC6gEGtBw++V1S
cUurDWq/EmXVfbImtCowos/HbtbCldm9AvhAHP8DCS/KsYHuqvW1owuRQh8r/thQ
NOn7KDR9NM6u7EygfvUlira70HI8IogCaWewN2P2xpx/JFbbQN5uPCCzZE++B13i
xWA8jPQWImL72sKCBxVeFU8WIRH2RxE/06HrWWkRC31O1mXsWk/xHUxDFEnCHJvc
N8bZ1W9539fmmkI0CJ93Kl+2NQPgs7yLj6r05gonsZKGXlIVmvJAPao6cSWyicqW
9WEFkOTwZzbavdXKReMhFPah20gdjRIqiOd7QU6Mjln7AztEtA1th1O4Z8y++wx7
KRVBvvvdcw+EvbazXF6nUfFvRsa+ZPhKuW/jbhAcdMR8UWOsb3h9KwMyvG5/jJQx
OtZuG3ehZhNH/UbToKgxZVI/oJcoxCDdN03NoRWJoegxDlU7LmdngrAY+0f1k8ur
Rf0vJ4rPWyLVZ/BaedCekETYF4br+jveler215eWegsqt5/pyQCZp4UaVgu9AW/s
8/2QYKtoigDieiXqiDzwPNKph3eHDtNYjHQ/WRy+AavpSYh35G07w1r4kSQdG3+9
IyapDM4O9Jm4jBq/brV2bnKZXHWMK16pR9Qzj06iLQO6yeoZ5lUNMDncrEpQeV+x
Vp8xr7cbjeNGJpYTuBHAJZC3kk1DyiXQXCD4YsGmsCt5YOcQpt0Kap7k58G4DxoM
XPsGaCTnonpnyD0gRTfgy0Bh2fNnGaEbECKdwPRVdcw47jAAwAwieZ9jZVkyx3uO
aNRFbxfa6UVVkNfEiPtSmNs/ZpDUGK7OgOV8YLmnWENJNCcl8I1O3R0CjYzlSVdR
qhWNo9BGsv9roLQAIVQdWwifLftfyhHsYKY1f4F3lgaJjTvAQ+RmPgz8Zbra57VE
IpBFfQXFV4Mmh7wG/35BVYSiiMYiuMzI8DskzoBSTQYodR1fKfpgJOs7ya35NmZc
XZ5C9x87la2oJNGg/Il3+nzeUMgPkWn7/TRDrAxWwTHWv4pGyuOicAEOmXqGOLtt
SirlMA/1365cxqiiKQ8Je0fokvtFdZSFkipM9Mo4EFMtdC2WTLEH05k2rFhwSR+Z
83zL301yFLBZBBBe8PPgFJcdsZDjs8b43pKZDOdXxvqoadplIm2YXoy4hAgHsWsL
9HQcZRpB24b971CiVarH4xqEWgwUdDvNpVXGYBi+6Bu/UeQH8EmIbHGOJz/wuAdN
H4vPh4NNhXKL9IBAGksvWD+nP9SJoi5KrQ/XWB2xZJVMOKa2E4MwXXfJtHtIbXXs
WctvTQKnwoMMt0uwApeuzXQMEs9h4ql5mXMoB8KzrzBW+DsmHXLrFa87ZawlWcKb
p4QB+oAMu771NK33MGDmUwEto9DEh0xLQjra7qv4qTACp2MUXGRHAaI2TAsHjbt5
GIpePLkaNcJB3qM6Nf7l5dgCae/Xf8bC2uU4sEfNWC1DuM/6sYbYyCJKxYbsnPeG
I4fkk0VCeVKJY/iGHEoX8PYhx0NJiTY5PIStdNnAth6wSCiEKHWDQtm9ggsfQ2r3
9XYhJyIsJrzXwBKwV8JOny03sqOY5y2j1q6brkyVCAqIZ3E6zSlNZzPvqjju034u
ZbFI/5/7Ga0S3BW+OpcbW4m1vqLJyx4tVnLrkSe7/ktoJGHFGz7w7GaoQHSm0KAU
cgYg3UZ3kvrAFagZlb8seLYDo2sRoVteCI8YPdIPVeYk6lCIOYHbo1Ge7Y95Gkdi
iJpjAx9hQ4ubf3hrEWjexBJvWZaRiX1/AD826F29QrYw9yWt0flWDlrTmmEIUzB6
2NChVqxEnNSONY05ql7kycOerD2I/yQwPC4+tCIDrBHWNJseX0d8wQFGcmJ6cJX2
+hjAJqJW1K+ueYrC4azpaLjhDspy2fjzp08jZWo1LnQXdFoMMvcYndYkmNeVgkFl
5TA0qGvPru8LnW88AZSwEYLyZyIpMTcRw3+TBPnitB8F/cRukul5dFhZFiTlJ6Eq
aogbdKEkuzi3gIKAYsFixyW3BA2BAmBOe/XvwdMeZlrQErmFRsNhCF+RcfoG89al
E1ak6j4QNZeaUrJSh49syaYBGj9rgemDEv9N3DHYiIGAuZLjuqO59FDRMTLVQJ4q
DjNBFagI2LTIppATg+tTf5VqTzKXsTNpwjqbP8ZeApnPB1t0QZkiqbFS9IP5f1om
suo0L5yAT9CfDGPWRYbL60te0FttGbQo+/ZkXupNMyf/GD64JDCmXwhYJhWonL+v
QOhYp0SqgguLNHAbKaq5AmroH8EYYoTSO1h/8OzkisZJkq6yve602keLlsH9ZGGD
M42LjvSpKFFuk5mAg6xakVwReWa4viy2lKtmGr/fS3/lhfuMBrBwRYm60ZQyf8Mr
tukNJp+lczYP7z7AuhbNYAnVaiKP3vtxp1j+1yiYJnEzJKhyVzE7X/bMHhKtRUtm
TZTzvnkXwatFOWZvpLYyGfwkedkfbF4Hc/yVWHVXx/jZC8mm02eNHjUZC4n4JKH8
2E/YkuFblYS5375Y/uMlySEV5lk9Xeicgt8mcYDufZavH32TLLA0ZNBbhTTv/kMU
K+moIFYRyWvc024biJ0CHl8EAxCc0XLxo7LPZKx/NZvdWdMPlWZtodEZCsVWl3vb
C5C1N7NSMPdPxS+KEATftNrguj0xD2kID5PoFWmu/A5OtGLFAnCO/IOND5LuY6fb
nKfJISc7fPDW+Org4RUgWTQ2WRkkfyE+h8Xv4uq4Y3MU18ocwa+C79frV4spKPWt
boNdosRq1Cj3Uf0af60JApI3RTrGCbUEpynoOrlicv5rnzp2u0j6f2s5ESxlNOTG
ra255a+tk2ZqxsEtdwrxce+N8I0ZD6X/3unLJ057PBQHrVn2jKNuwNRHIg1xKXJy
JTJrwXd8XCgGhlmM8amWkgI3OFnyNSR9SZZZOAq/VRmV3uZd46YTsJM1znt98tbJ
5oNrm7XIgfEgWeIHVOO/g8FJkKdPcX0+y+uPDtH/hZ1S8jMD/sTxhicr4L2+Obtk
iHjctOz6l38AW7cplh0lyZAw6HLQWFb/2TeIFniGx0MbzvZO7FwK6BErBelQLGX8
Xzx9vADTdAnFhcfx2+yNCZgs1WI4iBjYHomFF1bbgBAl4b3dw9ppbTJ/vcG4jcah
LcYqED/hH9XxHbXV0fj4UDkRzOK+jMYMakVYEN22wFt4hMCIMxkwgFNcj6Ru/+NV
bo7vs+FTW0if6kIceDoWBB5k4v6X78c2dPX1R89GaJeXODYMa1qfnrmuGTFofNIx
Z7zZGJcdLgeiHuyvUDArVCtXOolhKL3FHs4O/1AojszAppPZFIAWnq2eiHybqE2j
2Klf5+qw8VuraIibC8m02hTQyxELB0+tEICrQhmz44UYMs8wyUWjQE11Ids4xuvr
U2O27Lntj4nq7DuRtNQmYRojrZSSS0oeHJk9clTe0ossj2dnMpipBkkjeMRaCMTU
48hQcPjJ5YqLCSPqAULtpBH+9CJYn3O6hP11H0jkvQitIxQc3bi/QJ/5ICEctdUk
qD8QYMrJGpvAt8TU1RivivyPLOqI9vu7VOpmwzzNfNJd1j3SkNNHPArclwIijW1e
2XNzV4kwf1dafTHYLOtZxsW6JsG6pYIX9jtUT0Fq0MIAluPOKe7g6i8IU8cgFmZX
xCf5kECEt3S5VSvK7EvTq9aOYZehIMsFLYusYKxHvyjjokhtG1uHDig8lOwg7uuQ
o6YXq4ptFbQcnHlk+TDFBbCypu/PfslbGEikMXnLKq34OoDBE8Jm3WK6YegyTzYg
62xnlGq1PHno1M8bFrNf/66eOkYGe3mBKewGw8tuFQvOKR3h7X1rAdRzbv5NSzK4
NfmIitzjzjg4CucVw+IPqupJhrexkvBYPW58KpdoLS7eEl1XYlO8AcnCZ9y0ZSVE
DGQ/F3Uqrvy9mXUGzKcKPUWeD+9yys0lNPmLOZHE4xk/GcCnJ3kiWh1qwHkgY2f7
9SO90maNd5t5KptmW5iBP3vssl9b8OJ8tGJV8cFuLyy83G1W98N7C+8azJhMp/Kq
94Df5okq3peUMO7LBOtdg6b7P4WlTpSijO02glQLjHGiMbiwFKFwaMCkmtixmuh7
Pcik4v4zoyJG+rDlR3e48MCN8smUNj/si/c305cKSYvx6HP+wE+7RfowXUBp4e7z
mp0MWL0VNq8lpunR/NFvf6n18qohG0TIJRE8RE6MP4jvl5rJmo2s7U+XO5MHsAeu
uRisXxBErMcBlHsyViXEJEngKKI9IXqrrCYDszXELCSC6tv79bEBQP6azctVQBEB
YFxMifmCgUd/W12TTL+gcQHV2FDgtg8KztEDiO3Cxiv6INyPKWZUQRuojSEFY/L+
274wlH0rVWXVf7MWFWKIpZlKm8gl4+Ge+ctulLTwSM2fVPGmNqGdwORjjWn7KQI7
Z7oA35YpT2wCiChYuk9o9In179UZQrqLRTGXa6TqNBfM5KSr3MZjFa12cXhlK+2k
Yyss6uCXaKJfzL9Bv3qN7/Szex8faO8+TxyB4Dfa2t7UTX86IonS+H7G/Yq9NDOG
u8wshG6yWtkIlCtCoU4GM46ewPGSWNHw1d8SGwlaTcvktaPeRsDFolyrO0VXNW/O
mlC7KUoctnlzxe4/bf2+ryreO6gtK932+4eACwNLS/s+/8HVsrxynptT2CX8x7Nr
Qm8M/g5ug5im9CasizwFU2/bJmul9g5qZKIyyJsgmzq7olu6V3iDCF5nWuONqYbF
FK52Tl5oclovX/jUurAkdGM9mVOr2ia744b/nLoi+gJPYe+2w0tvX8CFz2bxpIwX
sOmPLptJeltqIuR8vmX8la3siNsrcTVwYxCaT2/OXh4N+BjgMRTWjBmgBWEdaQrZ
xTS3y0zDsGZ3GYJqgUwbQS/eiYXTmcSsX5QMO+x3QH3kiN/odGeEdLDAsfOZSCw4
IIApc/un/AngVMt+qxja/BKFEC9N2QZnjQc0eznbdMXtkpdlHkcb2nTeDM10fh5g
LfLn5Y1uBt67/+ERdzoXIx2t/so6LQocbaMi6g5l8V2EWWV4XrT2cmr1MR2yp1jT
UkIx8kbUn38SSV76vbHB/Rkbl7qAFutiIs69nXDEEDhlEllX2fpuzBFeL+jqOruR
xktXNYnXtS/D2zrlVaflv1Lh+IhTuzgFrYu0ageUqqWz/ymKnOyMN4RdEUjX4K1D
G+Wh6qomhw5JyxaM08I567sLIe2NWWVbUJRBU1sOuNO1HhZCUMAUfMLcfZup4nuz
/+b83xjWyprVpz84LzAgoM4wIaaNr9RwpQKs4jqGnTw3Iw9+p9APY8C7ZGoydDSr
QdF9tri0Frkue8tSxuuz5HpYhm6edQ4ZMc4NelRplN52xPHPnNkjDx57rEiyOHGt
DrNtdaizOCa0CRzy/ZJeppsELAQDN8LfolSH+jVg2Ff401lGVNE0C7JNUZ7gHCcV
czlBi5eJDifZAjTbAtduXQjq9fhPc6E+xAmTuBtc+KZ3hNdbfPBqf1lICQWPHmNo
PDDzjViIgQ9lPFDvAXjwvcR/KH/v+mThaa5EzjdPeBi8yFdVXI5GHzcGOy5B25Zk
kiR9IeWx4IaY1gP8r/5qpZC3Ld2rSj7ogCCHyHWLe5VlbLlmSRx0JEEaih978Uxj
92vr9a5nQ39KKzWvB1G4QaKkCGdCchHceuIo8vE4maQixAJjRyc8ZEqYciiQbGeZ
ZsQ5cXsynQAme5t9JVQKNbXpzmcjR8zTuaqLQmItTg9E8uju70ttcvUsS/iZf4p8
K/P8zrtI+Y0OlDDGoDVOA+eaLtjLY55OyJfnMEpSlR20QDIrt8QzfQBMYBtSk+9c
THya/u0rUX14ew4oLpEXWzgACK0I5QfQaQ9cRJUL77JTrKSPEdI1ycyz46H0YYIO
FOA5og+wSMP5BmQUIq+phP7z7vC8URkPA37RoyPolTqAMYLP+Ct4RA9F6C5Hgiyz
dJIIQXV1Oue6YkiOAzZOZQnkmCLrUyvel2+EfHjnPMTvOLYiYd6/DUN+zvlTca5B
dsmrcRTzeW9ZMWkTs+le0zBEH6OMXUCSLSCA7bzIu7nCc6PDc85Gn+25jzTWZrDK
0Gs4ulZpd/eZ+fUq21p85J/U5IKaWkZv1DMHN/IAGwGQwGOMGtiTTcq02BZMdxEu
2QtiM6/LxER3Ws71YykuTxeyenjhi2S/+/k7aK60gHjKavUfel4P05pQeW9t0vFB
122Re6zgZ80noE92Bb6u/pVzVhUEyV2eBzGOZNfWeGeTUD5mpBar6MLBZgPUZTda
M8/JkIU6Z62vL+jAW+e1g7VNCAfmkYjz5do1ePwIIuFAjFxMu/Dw4SI2NM0wJ220
/eIY+fQ3zUim9bOU0VJe6Tkgckx1Sj+2aW1m5lMl+FAW779zt9abBkZ/HzosU4LY
GAjobhIBpU/eq7zZEZVjWuv5eDQ78zszj9juA9Lm2N6FcirvqkjjZdDsNBwR7LFC
KAV2RZJRedutdhU1L4W0Z6JuSuHa4KV0xyn2C2tHFhipQzs6EDc3z9R5YuCGEZRp
Rw9aRU8Fh/i9TNxP3MqohWX/z04NIudcCe0hghEH8/A0p5ezVQJLEMmZZkE401oz
hWTl7av67JQAxygwHxwy/kY6pkequIqPg1yiVFZrxXn+Me3G6SuNUp45MwSasB6a
lJinQIdhoLrH0fnZ3zy08+Rw4TnVoR90MevNFCEa0ss1GRlJuHpdkjrMb3UcHShz
Wf/kRlYGVxR4lq91PqeMI9CSoVl2B5183Yd7/FiouFl5zNiHUek9bf2iYgN6sBV+
1zhpE9R1Qc0QVOH9zhd72iEGnYLxqOaAuOkWpb10Mn9fw0cfZDHoREScJ33MeUgq
IIr/xR5Z5mnVOmEQ0/oZnM+XDNw3idySzXKrtqLsSNdKkqcUkv0iaDZxldoY2Ipx
QpBKSEpYEiHUMGbL5ydoF/3oLmLJrLeSoi1rRVh7tv4qZGuAdT9tKbrAPLhr8MnV
QZ4GPTLJG71AzE6Z5L2pC3MSjEfLMxZs4wYIiWH0lsN01B0PMSJra2XU0Fjtz+jK
CqunXxI/s0TzwuSwBAQnVo/rfFd/avBJFBYmXTdCBZQPgsRfM7d+fziKauQO2390
IUqTIbdatJN7CrHNIJVZQSBiiMULFCCeRxnuvI8JJLGZuw8iIOKcJP6sL4iRxe0j
NYLTOckLhMxh4Lt7CiAJEYPNKtp0OQk9V55HYkvSlqQ5RmZbGr3ft6EyBucQxGqv
vbMH3R0m8RcED9PtWahLl0oMAjIprzMAJAyHP9CMfYFp7rMwJU0RQwFPRam1NPxA
HvQyrPwNODwn/NwUkqZ6SZ+JpKFj0yqf8nWxnNh8GXFDnL6t9XxWFIAYzf7HKppR
6/ye91sboIZCp9rOGSAupUI6jSp3UEM9+AnI1+q32hlCywQVouDyKHTsz1hQ3ZIv
8eXG5ZrmQAmNcVad4Hqx/aC3eCz7D+vXOwveZGh0Ioo1v1FKmS8J9gvCitbqz9l6
2z2+CrKWIO4ES4vKZ8n7dj6nHPselaHsuHo485ccvu6zyTP6YyxmrVPc8U0QaxRi
WjMTwZ+aZVpWkNDA9YQaAwoZiTDCzJeejqGAVoAkMgagXd1AFpCtce4dspOs3d6J
19Q27gYF1TxsA6E4MXmGNBGLibdyGE/dVkno31omh2kXuuSi3R4b8V918qiI1pbq
DYX6ZlnvfMjHk2z6UlwvVre8kVexNn0eBKU/24oHa5m1UPjyDkEo4FhVjatPml15
rg3O/zoTo1ToCqxIUX8OduMH8VgfQ2ctm9t6ppZXa/FJSj71n5GITh9vUa7g6AEP
bTsuBjVMSNPNXVZA75WAVcoAcbJoTPVGzlbd3iT9N/5lqsy3ALp0nB571PIZXhjZ
k1MbxW8rMQ9KCIyevnY9Cf6sJR5cGQqZ+fxPaYNGCnrvZSpikbjH2uFZGrOYYxrO
AlxpvZdJ1VewOuVDb/TGg7iXms9A74OYefDhDXzPhdBSuNhRAUhsognuWdZvh2Ym
En0MhJzTldVGZkulMQd5WqRywZ4Os9QOC9rAxsX8CiMfdj36JybY4cbH9BbBjHll
jnzIGciX0xEudshoGKjDUsylJzf/6JRw01x1uOVOuROgGY1cadRAIx2Q/uPfcDfN
dczL5t6v6TTVtucLCWX7V69dURNzG/NJvMad1UlpKo6lnVGwoG/gkPKTm6530V3m
vCrjrGfB4z4Q+4enegxUaeAyKb0gyLMmZSpqrRbUzKLo52WqWzOMfrmOTvZ9Oq5e
LSPosCamDzjr2gH6vPxP81T62qm4uEES9cdQ0faihytAbR7BtSUFVbzOarOA/jXV
kj/2+Juaqe+ZjftDGncXYovzUgJ6TUmsN3rzxwakolHiI1wgyp5rVlE85HQX287Z
6tbwMj/zZ3nqeZkwe/G9SCoCTKLIqhiml4tlMHldFS8K1mvh9YlcDZmbO2mK4C69
tBM++Y8SLUDi8W6UoCq5VTaF72Moe518ehRj2DDlcPI2r5qA0vbG/zRCVfKo0nNr
QjvW5q3tMaRkOdF8lga/i4H+k9cTC+JJ7/nIofGbN5wLuApOl5VEn8rcDW+Zu87e
MRtlZ9u7tNSMIcj+XNbUpYrKbu2phvo3fbWE3tNFLYgeWBP1//2LvoS3IeROnUwQ
8vrEQhtrxe4QLnPd6PMtdUlnYT8nTO5j+dMt3T2BBDcjJNGazCY9HKF7hrwOdKYx
m1W2w2F3yMQFlx9o0sA+I+RL0Mdhi1kuGnPPTwXREqZ3ts7dwiuREbYHUd+BqGid
rwsOcxgPmEV7SOQvEUgqRWlEPyeyruoj8xLynhL5kl7oUnfu03KzfQu5L934w+yp
Ah3lp8KRoN8aHgjjpVLaXWv0XiC+iGCPVl27BpG6qN+hXg6ru3MzBrznDb+qv/Ye
7kMJz+nZ1UlxhK4SJHTrMh9bzeZ8B2dopo7zKYwyJJznnBtlxxF2y+5QsDTM7TJp
/cy4E1xpHFlouMBPSGQpucR2aUSvgHhiyNydb9WwWexsPKN37q3k2YnYEvkeEIy/
fIWed09ENKc/d7ZkDvOpN/q0u1NhrainGMjkNW+pNC52JALvj2pZELRfmysMbCnG
buSS0OtcodIwEOYZPWwM4+fe90XZmOH7gd+5mO9bcViilHtpJJftsyUOrd5Ddy+5
WaZLayhRVTG1QOPa2D+RjL9Z3NBtczKMspttWhuJROoZJ7miUjtCnH+9Wm2pTS5Z
IYwFQbHndcDuwGmqM/ZZdSKfIVhxwHxhceFSOVG7bM53Gxpb/msfSmRZp4ljnwZJ
joYWW8Sp4WD8o/mkDq/+cpxtgOvONMKPBCISbeNZESvktIE8H8rZAMPWsHgZgVmv
faw2chc0R4vI3/Wg3HO7cjcNercacgYB/kpn3XTZdie2JElbdlcTU30P5rAYXaBo
OuMXabKW/iUTjdk4SZMEcB0I1l6f748YG2618i70oeScZtmU6OD1o0VYVUCpQG3z
YWWX9aSeZBVgDxuUlnSgUpc+XDxGovgEdsCTNQD7OwIpoqE1+034G1IDwSSY9TID
TPz1pMR1b+3xWf4c+wrzg/HYusqy5wVZ5bGwDAqTYxEtX3WBzAmxgFF2bimfemDS
1WRCYR60vBwGdeIYt23W4KjeiSy9Te6UHN98cQp81NWsgtObG72Z6gJoLbK4YZWc
4ZktJW4a5lGXqdjQXnZgHZ4Ea1aWXDN54oxn8O64T2nNcTLEz+rNO/vitFR+tLXO
Zw7gSH2HjwUdOyFRMah5d3wq+0BngGJ+kz57sQffoarK2mpjJb0WmSG1aTguYpfE
4TmPa97lve0oq26pkSIuaNv99N1ZfVdrjne0Ri9BLDasp/5e5RTCeEGl/nDb6E8D
1lsTSumUx/kZ1/OvitFnLhMeA/VtT3FskVOJVdFTe7oYtakgJo+1AAKp8MQWk/iN
+4fbS+EVVJ9B0uE6SdNjPnhiMjFIGm/UXgjv5lnmoEwgadqbOdPUdVjdcmxwGBC0
w2C6ufVSeEQ/noaQaUVO5r3DGod1T3Ez8BMK4aKYGJjs5n7Te7pHBgIASlQp0c+/
4OSEOBxLIP/ePh7EuX9+R5FeUSwvlDR2bh14Fs17wQPSI2n4mk7h6w1dhyIBh53x
NE39jcFFcyeBbZ3TgUxO/gxmourrxg9fjjf5cntjWVtTNz52bNTcqjzzI8Cuj5+2
UXlL+vF5hBoRHL5C6/+silisrzlwrn12VlQ1YYcvTcqn+fooKybSTYorskRB+BsJ
/HfCW9SrTL4WATJHm7jtZS3qhv2BDR+vM/blFFrXdFG08SdrsxrMDNQRZZ8g5aKK
S/NxAlT/yKD2aoAVp/D6Nq4WwrGzyo61z+VZCYPEvcG80OrJuP2Wfun1w/m7n6mV
Jn3P1KIcGmdEFoM3pJK4mxPL+iiAvmD63ycKndzLXfEN451UCLwRUq4sv3zeNv/C
AXvhvNNN54SYAV/EIvgfd8vgJuPCXzgp8EzGma3MJNlTB7aZE6+vF4Ca8+tb7Ewr
Y14DkDKgtqy9K7d5YoDj0dyaPmhnvIkdcEUsTvihmakoNMMwIELKpJ0CERRAaXUl
ZGBTl/Itq9wQyBeVE2ltNx1tpqRwtzh0QY349KwheJFUdlKe9Kw3sKIG7TfPvJxC
xYhLfcDPZBmRZbVpyJvNb5cHFBN9DRrMyLSqPgemx4ZWRb9KTZHoZnBIEctxHyKm
xRQMx6arsG7dVsEJkx9iGjThxq/0NJ6bYpswKA/GzhJaJYrKwo/6CDW2HIVCnsvc
Ehtx9MEaVqbqoyLotj5/IBLsymhIobcy9/5WwnZvA0rAPWfIhM3xVf0LjERfRSsf
hb/oiprNdmKJlxCOfe85SmFG2OiiE+BkkiMlq28ALk1jaFs/4SqzfLtpkR2A+nVN
r5zi2WxFwO8O5G7X+K29FgjEktrjvx8jwBwevRu9N5RGl/ZNMn/SjdOOGOqug2GP
aoL6d7CTAIaSXZr+aU5B+c3D3t2ccqJvK1PuZBWH0Hbk72AtqkPGZ+kgRHpx/yJ4
zb21PeOVPIFhxENsQ0j59ZubM+zyVmmn4O5izTpERv8e6l2+gK2iKzfy9YTOC26N
m6s7K9bUyTfPQf4VZESKbsWMUiWEsjVp73FuQKqNdcORQ/xsGXO688QsLBJTJZx+
Np3qYz9RqInATuN49fbNXsUsxhL0OY46SnyY+5g4Rqnbtsq1PcdLgsol83RvScsi
7THGMEHxyegQD0ZlmTdDkmNgih0LHT5xxb5oWe4yR1xKv0gDfMQzzqSBQME2Fx13
Iq83wkxf1Uop8vlMvbPkDovJhgeV6w+doEgu7zwoHoXALkJbaPV5DMfLnXRNQ7gW
oEixfQRVpK9xlvYhf9Z0rZSGraUiIzP5H+F9eDK3a9HdRvMQV7phAc3raH2MI/r9
uBE+b1ur1EHL3ZcqDyqGuzC2gYSiklMqJBhpq9uOfoVKrUPAvDY2ysSHXtwasWRO
yFROjc+Ygqr1gHlJhWMoJvq1ksCNOPeydFzldbBLC13NsdNfwRsSw08Jpr7TOAuM
cjxQRxJ9NrsoRlDB36dJaWyfuzSe7TKUoOzNvm9ZSGQaftdU6I5S9IIuftz0v8ab
XiLqWnpfN5gr/Uhxq0VpBrJfeZ5DH1tuTquy9F1c9GUmvvjKWYszrW450yaYwmQK
Tkyek9nvvVDEJSYO+RpiHCFr7DY//EuvHr8QSYn4u03qyF1ftNwAoy8NLXjTcd7Y
uM8B4Hdh9E8xC6lsyTIOR/X0MtDreTeC50PjSpI/LPj0dKKchXxxNNvpJ0y2D2Md
zd2+O69GIcrexWhR4/TJK8qw66LrC59nnNsao+Akh9OEMQwE8yGC/YKyR4nSIpZk
fFauQVmP5yamTJ2148228g6sNX8iXjDAu0q2NkfTaAbaXjCLORxR+zdtAoyyXZHe
W28dXsIAQcmRLPoc/BMMn0z92ZkHsVQLchma6jkqM0KVd+euxI42LZ7ZjyXSuWW+
U7DwBGoHTuQjJgJAqJG5NTmseAU2ph6goJcTBHLd4lMW7K6AgrgxBynhH2mrzePf
qtBdNAk0+1xLSq85x4146Z9fRNKCkl8l1Z8CvWk/XALj4pUTnsaHscVp0gwmBKtN
aYXBHe5tndL/d/p1utuXRdzNIXS3PnNIiczW9hKcbDi/CmWdGm+gzZWRBUYYYWhc
EvSMYKSI1cJ0MOSrCnUJYGIf64Vw2CjxQXAFQnuf75lmye8JOKymkRrUFZmqJfY3
cwBSn2q8fbgy+k501bOA0mZgEZDZnbOcA381VR+C4GZYGsDaWD9F8l+/JXF3/0c8
Px8k21rOy/4M1Wd41cqFMdgCAN5N4p4SI9M6bX8+tSyOyKjfe3IvcsksOdk9+7/r
fQS6sx0OhR8EJk37qXv/HBomIaRGbvPpIHqs9x1l3Do11fU5jLMlsNCLde8+GkuU
bvpxhZWiOn3qCvmvAF5v/uZhFRug683VpuW3km+T4ZOIWfSp5QYybGtHqMtQ1ozO
m7VRC+/6umz6Qd9CaN4IwXG8yYz56pSiVgE0eb13UMXIi0HdeRPmd+EnvYkWNv1s
jt/itTXrpaHZtMExLHXqRqPZ4GKYlke4NGWRcDsimM+kO+IqF4VnsB2qM0Tdw9wg
/S/ltWiAgIctXdVI2ePH7+8lJpsVeVPapt+YIhs5QFVFrcwCmVBktJQlLWilPzF2
CsO00hxuN9S/w/rSyzf2tLXsMlgINh7gBcGvTnZ1uxqLgx995Fi5GxVI7a2wsvVH
puJTZ5whfXtQuewI3QDULo+F0jOUsabkDsvRPcOlcJZxdEaPdxbTQ05hc9UhqiUK
6fotctlqBF1uvPf/MbZdqb+oHXNO8CLjD6VxGwPCQAVaSwTU4cxCfdtZ9hjxsZMy
rJrMxLQFROw92AvS/L1IyEFahKshS0eOYbv1Xii8UKcNqSOl4N6mFUXFPTs2qPN7
uHM54hSqyWnJsm7V1B0vzDuFQtSvjLW7gIwpOFNR1TtcEo4ZyguBns1kTD/ycCQJ
hQrMdSbJkq/8u2cjSZQF/1VaBG36FRfirGxq6btE62Jo7UnNY0fPS8Zwq0jW9UlJ
q6w4wpOp88lQtgL7uKxybKOtGs8IpQqds2wgdZePY12/IecNyNAUjHrK+P1f45ja
sGE1fnT8zr2KFh6CYSym7Bn1mBb5XWz/xXNPdBuCFP8QTUV2831d47I/E0pcAFc5
42tSBZBPlZZ6b/tPyb5QCAraZpizUvw1mMGkqCm9cLnybtQD1zG0zWEyztCBEjIU
Kxxsfox7sDreRS3BQMpp7I7zKINObC3ygwRcbWa0rOSToWv42Uf+e/A8p3376nYX
hdnuwKxgnO5AKZh62i2CLa/+kl/OHZSW6OCgWyZ/SkVLNNN8pQ8aMdnCCK53qijM
vRGoKylUcnSHLrR5pMzDbOFhXfHzT+knssXh79BNUQqRVTJneGUYpRMMoDIgFsoC
zTnj0t4Y7v2f6dgSitrfvRMzsvNFMIrltLMM/Fwz5pvtdsFkXhusChTHJWK+3UCA
sRnNRxRCvm/6Lx9YWHVJau/SHN6NLzgmRGJh8a7FDF5KCNU7mR5JFhuEhmrhXtNi
gqGoK1M4imp0APj/RXGVh6OHkUjFjj+s397MkcAwROXSciUoWE3BdYnGxfA3ZBeK
ERNTudbEE+PVXYzOWe+DOeB2ZPQTnaqV2SdV6OI0xbFkDx1czQjfL6kxgE04mmJb
sxrQQ4wS4g0ht1oIQCpaspS98bgIbYg/W0Py8wMF6tTVf/d1cJpVMfs6t4l4DihS
eCdeTXS0cVhUkWv3JOHEHDPW3sZ24K7XxhusP1bqAZdKEzDc9mcydV3+sm5LwXBm
7F8XTkZ42PRpp2fbGxQEADpFH3vZKAI+8A+hg5fDM7wA3+igO+IK1cT5MVpt0XfC
EdvISK45bBVMcf4ocxrhkunVktRryGqfCzW5Ld8EUi4GBDbHpxZjYvoWIhFcOVMc
InxOUn1PIJjh/2Briu9YPz6IoEkYt6vWJapyfkdWbNfQWdPPhLKovPM6lZ+5X7p/
zJXZG1gRVXOULiHC1izDLXuxojs2O2CvBSlEnA9FsAdIIyZUw/yqSisvQPJ87EYF
SvrxgmNLFCELPA98OZYS0TQ+Nrm3zox1VmwFCqG/2W5cSLaqaAJnLuqkOrZCWB4E
ipPOqKVfJ+LnmiCFEwrr2frkxqtu0xrcRPLsQzm7GkZmg8gCiTv+4SAQOfMPTlF8
GVc4IOTAwzocBjdJ5/5UUEsMfwleKHEPgH3AmHt1IpWutLVT5Rfj2oXwyqzgGujp
esG5/qXUujW0gWq//kFaPrTjOA7kUXCze+9XT53Rvm+F+/njmI/ahaAadrkad2fi
qB4q+Hbu6/AY1X9tqh42V8T8Ecc986rxp0DNKm5FXBjpb5bXLgcTIr+e5gooAGCQ
sUXi/Wx+RUhyjCyw2PSIkmSkpe1AqbOLc7a3G6l6Itw4IOb75l/g46bt4chz07aj
dA+5CubcLKzZC5N8BjIqyXTtDKb28uqcJ2iVg+B/xo87GqzuLOJLbQyFSC0RuIJu
pw/eygtQfi7UB/J9SGBiBMhwBN2XipSc9sgJzg1w406aI4uJtd56eupJFJ/9Cq82
aqhyqkjqBxjE2hbPLUuzp1XuXlOa4WBNVrvvYAaQ4xvqAbtsKGJNODkTUezlP4Mf
meOzvblufVkyyyvjVCvsGJAAHd2TPKuhW7aZm2CLgSG+4dKfO+gA3zMlj2MJQipS
JLlVGX6ZdgYvFJ84JVsV6Hq+9YUbgq6+hx9ziKnwBJs9pKp/zgzvbOY/BOoSRKmE
Bb7SsyL/cluJ3gCS59Sz4XsnJPullMETW4GMrgJ6XP9vQrGj+JFS95BA2gXyWc0/
6P4Dt7yTys60iP/gzd/AtV5WTSaUkLPB4tPx9zkExA2sp90RfcT3c069YptOnUXf
ot115s1+vBkXyFhzEAFN69iPQu26PvKk4yuSJERJsq00vZiKt30ne2+8bNkv6BFw
kMdf6SeGpHEamXy4UHKVOnkEOuuLTh1x+kiHIubVAcE0jOG67lRtGJeUS+TpVedA
zZlljN83r6gjRsofYibjePgKrfwzX2GYJlFZOgyzkFhBLHtdgwmIPZdjNzDp2f0/
whdLnAZfBE6lS3JM9MiTEbE+J+NvfsIQQUQJJynx6Mmm0wpwz98nGwF4LA1xoL9U
yNk+kqYqFsZZabuA++ME5XATqIPeIEzkXxhi+Vhl7q8DIQiG3nItEBkjHqARoRVV
o2BmDPA9epfZE/FZju4Fe59gfM3iekHQJWZW0j0RLSkFRi6elbOFECHc++4a3gmH
TZPWoQJx+CiruAg37SXsbyg1IxhLfiTm8MzxwuQEngtmjZm14XujHG4eGt2knDi/
waCAvo+MrD/DnFQnU0UtdAUddvrnH5mgXcuJEQDwhRENFdbCBFORoLR/tR2Dw5Tt
2wqTLvZJfrdEpYy1WoSPXQhfmKwlFcei6YhtT4Wu3ciwde9yU1Bat4fu+QfeRQgQ
RCPJnOLL2IJyWBxgD0Ps72A1sNEfcGyIk07lp6NZTiBQulmxiKgKEj6co1TGPphu
YPwncIESEJ6x7OPlkOr7lbyT0b2x5cCYV41QPDq7Uf6l3s9hh+Bp7EoxnxH+IjkL
8iHWk/S0hVvzYgXpG68iSwio31Mi+NEsmuCssv1mjTr3ISoU5uTtaoezmEHlqKo2
aIf3Cd6cvMAL+iBEc5dyBvcz/4bUKAJQ4mWa0RplGozsrPpteX7mQtBN+CEakQEZ
DHPSZlupv/bMF/NkbwcCKYIRzupdlWPMLZGBwW9EDwLh5FJDO76mZpWJCFJTY9JH
w1bwfqi1+m3o2lSJTNRbzdfecg1DQVh9+hmB6l9lyzD8KIxIo9/REvx/xDIiSQaO
+zpbd72WZ7tHUYaHJD9xYgMD51mPu5WW6oKCMixTf/pjfW1cG6C2EGnfIwgDJtqF
ZErZwB4JlCS8KsHVDvEgrhjn4L+BC7MzVDxfI7rENfYMVpCFj1zXiEPE0O5fgUsN
3cfe7JeEbKM/GFrI8U/4aPnfv5bvzw9m29sYDATuG0qe3uUWaXKhzKFDps4aSa18
o/f/clPFtdtnpMH7/AEkI+tcZO5cnvoALo/NMLZMS9ggfOaYrsNr+3nizclNtZoS
Ei35odZTQ50OoUpqM72SXFIjQd/HhVU3uCPM6fubqj1SA2O6o7pQvsr9iCrXQQiy
8HahDBNfsC+Bog+WniONhzjAz0CZzB4IW8so36Tdg9R11WJQvKgBH2J9qnlWpF8y
jSDzITM0YwSzGaFMrzmRTpHHBvWwQQOdgGwZHNY86WbCgedqZO+SZ30Uo3ps6wQT
84Zc14c9jnE0UyOpkk+zs43YIwpvr1C+fS2cKGF/Euu9yT0WA9QmmC9QV00vIyaM
ZhWgtJr4w/jIZlqcDfQQTw4h5cdPdE7aWHjBc4L+aMLrHNC38ZNUtdtpapjy3anZ
+vExAOTtr2OYwhNzkN78dbyC5le2iwclAZIoOVooru3xClJkAErb+QrIUVs1S7St
Lojr5FfbYVwKLq0TRMM/8yOLQY7+EG4zhQvcWGzsOCmDvTyYv9dErKYyW7GZ9ApF
ZTL79KvIW9BtMvBI/H95fmkE9gZwo0ZJCMitxA3R0SFe4Q5LCCPy/SPRH5EuC0KT
q5ypOH65jdKiQE6JPOtlaLAsD3v2RXUfJVPW/qPzTTLZehYJ4k5dUZXAsRuYBPsi
I/+TJjnUBsA+SVtyqU9T3ZjCqJ6P29LWmC4l669KDlEIJj0BYDQ2T8jUTpjCdBqw
YvxP0EK/qSxZzbPiHLB0cbW3t/auvTD04ucQTuFYT78YrRAbsB5xobfkqcr7+9aC
zwTxkCivFU/bI+liAP8qs9Pi4ZSF7AdyTjGzz+0yr8ZbfQL88eq0Pgmia4jOh4fC
ARYrtIGjXB8ClH5HBZk/MsIGA0cv/5m5oEWviyM3bmFpTQ6nu1gSoUFWUQnIzXNF
tQU05e3W/1FpmBR4Aepm2Fdm2CQP2y5n07IPvUKLwLg/9TEB2uKu8o82DPZfcc/a
G/8X5lTBrDp+ABZ9mz+pQ2YFid1lcuvipZqw92KwotnKe5KujqjXNs/viPea7JDf
Oqrv2oU5jFlZoyirTA4OTwxzkMP+5JmkS4mHJfnSdzNL+W5vSFOyLp18oRLqQ8hz
XguR/oLVbLsXaKxGaa2gYdVqiawvDcCYPeCojq29dXJ+gVaj9USDWtQlLQWJSXHC
wGgzVTq5D+/GQiG29Q2+LesUrVCrXpOXtW3TS+xOHdbXxQ9D+N8xaeLQ/cOuV04N
ZHGDz9u8cU3WZ5hyw1KTHEiGXsGDwtvhKy9OuPqqyizk47Psnn/njWJm9eIF3ta3
SADMLjKuC8hORnoWu0v2t85Yi5SKNzd3fE8UHmpWkc9WdMTiUUiWIUs1YC7/umyc
Qq8wuGH3xPzDGlxzeQEqobAyflhBTLZ/Mh0pRYQmz1MespL34eJCDY+TgvJNbvYq
TjVGkbHmvMYlL2Q8wEeSLI9WX2Up75dagj30DH8pbVY+aJ8HseYdDdE5OBJT+hN/
BCLZJaj0JtMxU46R6yzJdT27aij2YtqceEKGozPu9cgRE4MqpD9fgBVQXjhojuZz
pjvnNptWOm6WPPbpx9rtNjVBYtneVTLk3WQhPeoVJ4E8zAoi3EHi13Msm3p3o0cA
wXGkTTx2YiyGJCcL7LDfzRnTEVpFmLaOA+BD3G5mJxBSeGxgvJO59AcpvtgEv0kz
vNTc8RFhtZxQ72GVc2PMRB3e/0udQRqyalfRshEWXAXN8lNjLtgk/dC9tLjRNRWF
HOlW5pndaHYYz3yV4eO5AoS/k5V2EKi8TyWU5G2a/nicN2SZFZiKgzihD/PVURBh
F6RNZ75IZskdypHUjDsjJbySgy0MTvs797UPxhm9z46IJaFquyYfJLZbCXMFqneR
fgbFVeZPShB4raZ9dszjTDm4vxaGx8WqpbgZeGukR/tZaUTdkTBOIuNjo9dDx+P7
UUzdLgBnqEY4iYb+ZrT33qr8niwlVpACV9zLcTVadvqamSFbKFZSONcjb84IbvyU
TXJZ/2OPkD8IgSHiZej6gTTYxj4HAD80H1Cv2/T7fdhIhx2YAxcmDVmPJKYIXLFr
79bVrIFuahqww3m87vZUaVF3TvOb2mBEtyJ6zAItc4TbltYDvT6YYsfNTtQkaExu
0jg53QknF8tGeRdg9njG+ZZM4cx2BN6OnFKf4xIPaigadmEnQzDs3EINayLsCb7G
/sOmgFrw6u1tDRFylqHfRbnCvtEIcHhC3ot9laZQ74PQPAgYbA5J/E5R++qZgFzQ
CuWemrH9AxQztH7RE2LyJytZPexK7gTmaEvdugkPrtKqNrin8qA2p0a+SrhV/nUS
y8d9FWNC0OcasDP65vjq9ux6PSDvwKNKkuPzC916Q9PjJO46eEPkSRlruTBGsiD6
HqjalzRQQanFdYu0LhPesEpWPnxyociXngvdXYwod+4gmhA19MNl699A8d/epdq/
KV3PRwsPYoZGuhLLBEwH2TgO/pUnEiAJFIU2pLp0EoDw1BgaMI3JKKsYsOI00Z0R
c+9whLFbSekcCNhSBYWUUcCTV/WVzQmI1m5kWLOBrYllH7g/gQR1Jtmex25+cB3x
u9imE8vUQ0wz/EqCtlckdI6mypScCdvRZ9ziydchOjGtxGqlWTB80DVMvVy+PFs/
7axTmFggmeWv2E0RMs1rTbqcfWQcAF0rq/HbErqZobO542qB/h/9s2KjAC08wfPY
ZCrAQvZsc6v2y/HIdnH4ZdKPRP290ycqDGTlYhLO+z+Tki+mjQzdcnM2ZcX6dgK4
TG0L/jEd+PXJkg7duA5cC0f+0Irrf8gGzJRqYJF56J2PaFgV/AuksNvJlRehQT2V
fQl8iDvygwebBYkFFP5JqFd/GjNfGN4HCF8xjUKttFZ9lleT+iBgShnrnegUOc5A
D9ZTPOIqpA+jgINPPhE5H4Zv69TOiqsLwSztp6jeC3Aprmge6AOtmj1N3rYMuZQ2
M1j7pUrAPY9bZkz/ECg+qj/DIsyd7rczS+I3JY6zCf9+qQX1sK/yU2+nFoCyY26+
7v1ylhZ8VJBxLgcmw5NldQdCz9Qj0eefZATXSqsuM9j0D5DCkovEw04wvSvNFaEI
3m3fqQuIBXnGF7XIC7x/OlHVOyzQnOQ2ncI3vCug4kXYIFDZJ3h9Soh6Y+RVsIqC
Ws2lHCZx7sgqpI9sr87MPc4j0fof0icGjf60/LkyxPSJhQI5MLJ1vsxBohvsy4SD
HWcOAamK2jylDjJeAlw1cO+CABS7EivzRGmEMpYUi2dEXdw7wl6tNc/G0hdUxwTU
u4XpW4sE8q5FiEdLRqzBR110sUpP19mZ6XY1FpRLywnMM/RrdAwTORys4TyBSI86
MLlKxCdvYzawQUVy2nbPYByXe0K30UEos5elLZ9s7glpGQKsU0sIjPzz9lJcVHwQ
GJQ71KVAVDjaJn65QlO0sxQK59KmknfizrRX4b/4u1bwHwNZ6ab659Au1um2G0nU
FX50jrenoPYsHiGpDzSxZwKCx4uHi4fSsCcgHGUSqoa/0RiWKeE6HWDVnKNvS0Sg
Q3Q8/VYpQgEeW1q9wRW54Sb4QaonAhQuv+qVyFnGbjBkdo3KqkmH7pQEVuEu/oqg
26x5s/gAVMn4RFxp3GFYaB/s7Aj/CuoQIcoyDLFgKwLZe87XUHGGv7zL3Ofbv9JK
T72/jd8kI78IkAnnMpkdVW1u3yi5+UdmTl/1DR1odYTJMWsbArMJ5j1usAMR/Jza
5MpLtF3RBfgAP8pe46xGkpNDybpZ/1WGzxsX20tZgA9dT3DV2tk0sG4dtCVE0/Lk
3cXQ+evoDu9tQI4hoWjLQwJhizKGMHBUoDZ5t+0r8BYETylBwS/czU4hRfl4Eoto
kB7cIAZx9SZZ7YZAdks5rDGzsudww2ADp3qATbaXrVE+oL6i6wok3G6FyIaxux0t
ifNHQcuDYZVir56Dmf4xaNY8l2syL50ubY71+8fJ958l/UfFoO7WfBeL8+igi/uk
xcW7Wjd4Je316jzJyLVKtEc+kgLzInbe+CqKjRB933dasDbpj7z5Kb21HfGjCa9s
BBaoyPT1ztndhheVYop2tvSdho9HLMoc+20Qbg2+AVLPiQ649c62HLZYaBlTDB96
7idW8VX0qpDSaQlT51YFhhysxk+LEStTM65u+5NBGfbrKuKpK3Y5iwdlbdN24aJS
erMljEWAtMaM1RJHCG6AULMUu6nS7fpbFxA+vM/Bm3Zos3ymzOaNfUjFMg4++iYq
9WM9qIA26MjS82JJPp89jX1U837aUv3o8WCHl/U+yRJ3pFevmr0IDaCSehw0vlEH
tb1/DhtWdn5McDr7xIduWJxTxvSFmWqiRg0/PaP8jnGK13o109cYoBhvnEiGoq7F
/mZPgxZ8geus0qJde62UuFbDbJEUv/F6z9xic71hyMK96OkKA6eYfWEBtY830vgI
/MJeeOXYoc1Av+h2avkqdeDei9HBa48EW6cV5BZbz82tIKiR0Qd6nquGIr2RwdIr
Mcjg1gcW6bOhO2UuSv3frRFmzDFrrWjsoy5hStiGaJRtn47Yc1EmlENTovyzmNZ3
cZIfkh9OuE0wf5GJHFAVcOT93FS5q4Y+t4dfR2AEizwbt0AllF+GIyfok0yx/2iq
FllXqSdoNJlEr9BAUnbglFf1ke1zdTtbBbQAm8LeE2ir3XKU8NcNtmpWg8VkgSc5
V4LOVBLZQchYy6YMDdPTalmEXoCrj1vbQvSVFHWTtq6VNYuPOahUyji120mMuXh+
kmdcP7Wg/TyEs67up/yA1NgaufA1TnSojqtACIaDi6orIT8OIibaj1/8edJ+fLET
Aw2Ks0IJXwHn1//wH4u7jkmynoj12LwH7Jy3Hds1Nse+1nn+IbCDSliKb2Hs1Tid
ODDv5bQWymlg8ZPCEm2zsLIhJkqXr+HnBHkPotncGdAHi+DLh9vO8rbT+/whuMWF
9j68zN1aXKdSIrKc1ofrMC+Q48yxOMnYc+tSPvHQMcAEoZIPxb/KLJHXVwrKw5V2
iv7g5qCwOSeSLmWRdJQ9YzYS0szreJPUPHC5yd+YMAUrdiUPcgYy1Vb6EuDj+VVF
3nXawb4WaOcHYC2ht8QVLoVkoLJXcdA57mH/9yNmK0FA4FqbJALISmVw6nQNi/Js
XwW4tLG0s61nmhJnxILtuLzAT2zKnRtR8AUQOksF+E9AqjlY1s/nsRJxCced7DEP
85jqp7eM9yASONylqkYWuOG9/Ik7sqmZiI5KOttyk/63GQiAvBVVeU1ODt6Xx842
QpL5MvTMt0erzHZhh6v7gyKpoApdlJXzAG2ak3Z1uBXjdlGWn0emKq51oq9tlR0o
wJDYf6LTP/l9tJbrJKdE0exEEeaFL81jFbh4GT4UHK1tFcps+5zhkd8xYEZrQ34D
yLT8uC4YYFXKHG4wdRVHXmamvTNw7yrdcLIt33LQxJmh4v3Mu3yehFW0eGIllmJz
9jAMRYHYUZsBBZh+f+/1vSLzGTk68boVUl7ONhvVOmLLpWpVmRZ8mFhX8BxFhHof
ow+PQKm0GGAx55P4+n18t0npjo+l63BACA1vfPigBSAlP/Vofk7pj4tJ3+FA7HfC
lQQiYcJMJTcu/3op9DsWPdfSAcv+KB/GU7Zj6MeGoZ3qFKQQHOTMAL5AE7WtBy8d
9xAc/iri28BDhjh0B8iK4tLmHWLRVPbQ7U7MFI6Cw2IGpUwHUbH+Y5WdXpT/wE30
Vib9GCpelg2xFd3Du3pe+rOB50vin2LjC1QbuxJAU2mkvqn2eGGGQ+0ouVk2DwEL
kh3bXE3AYIOeJgIg5/KrzO1b1aloUq4c5MLLKyeE5mK46ZObQw4gOggNCPIuYvnk
iuNj+7RCds0iwgBa2JDkcZSfYjg74ltwFbmxzG8GZ3PYTSt0rxSLVNPqxltFkUQR
UZdSf6kbh93kqq2+K3Wi/RbM1168sr47T6mEqMiao3Tf90N2/38k1xt26xJ3WcSD
fwcClZCOk3XWMizurWC06Mb1PnKUY1xhu3Bsr7PO0FqwFELxIIEBoTEd46D0rYVC
bnSO9EG6RLEH3I1fbYgNyBlBHoVQJraXHBgb4Kmjz97p8TPFtjILNsLQuOTjKCuU
WeoBJrc7vOc8NBCNf6hoZVuheBRboxPr2iSlWMf2k6mMup1YsfLKjvXZnjpgQxSN
Yb4EEnuFW+Ffxa68slCLb62M922frJ3ewMVpOJmS3dRG8c8SUYTpBvq0opnV1a4v
Nc+8FKMnobEco5TiVasPgjtzL6L8mGAhXHq02yQAADEqx7aOnasj9btpaJabnxhS
sUdy2/hZkOe09+iczuTv/5MKcxMrqCy9XAOE429bLajJQ4wJB5wh7wt0tLq+ZfRp
1Jh2QNDSYoqDln9WLn8Q0HW3l7/o+HuVZTdSyObzMcl5a6xHTwabBShTPcwtc3wF
4I0OtbW5sIGlfLIghLNC6VfGLjMAef5hS/kmHyc++NhSrkbJO3UOzSk/g6aIpsvi
0nBiNjlxjZUZ7+vErhN1WFkUV/W+0VqNsamqfzgHAUwX5U3q2+9ruuTbnIdbpnfA
XpQsuc+OtWnkCWMBUw2arnNw3i1x00Xyj6ObueJqJvtKGg4bt4ERJbGMAQRt5LBu
1Uwlzv1BKz73Rk/dIukhGuB7wW0ufesZLDfomDfoHdQ31JPZQM/PlzQo57v1qYfd
4VsDod5faJnrOcInNBXuKeLauwQhMj/B/lpqGKkEIoQcDa8dkO5shgOyapOmNeJt
a2VdPe7cpR9nRZHIzcLLIiWEhGKwP3DIqCP7w6KZOsjLjaXFW1XeTUfAsEQj6B1h
psZV1XeToH4TIzPMZi+yGOPlTiy9gvLxVFbYHX5Bi2+R14sKAFXatcXU0GkPxhu+
58r1g4+RvBWoZvfDqhY+NzfeEa0Mr34f1CyCT+2Ea0LZhwOeOvfN9nqol1470LP1
jtlcK0muC3GRA0Zdxf5K54KnAp0Fjuen13TsURJa1C7Ij2eWbwOTRr+Xa/0A/TVb
oXSfd6TXuHLPzTj3yCqnOHWHd2UwpEAzNf7kuvzcIzksm2F2B5FropWbAvhOSTxF
tQyxKbUfSvV3QZpquaZjlaFTpyuKw3AHyrW8e40sYrEMXTGnd68TTK//JUeDpQDM
WejDwzpP+6ewNQu8Mh4CPrtYx4LCiWhwvG4K2aBMlvC4fSKY+B9bUercVU7NJY0Z
rHwns9vJx9v6fl32q1LRryLmcNZRDnWwszT6+P8z0gHi9Gn4Qy5LtF7dLSlJn8kA
B5iBz4oGoPozKnmYaMy6QXHmJtVUntu2BXBqfZbofn66zY2IwYtNFIZA5XT1DNLb
Ir6LifiyBMXoyisE50ofTnhBN5vQ++NJkRJgp7q3+1jLZH/uwZr54x5aMffL7SmL
qCU3a7UW6lRqQ4/xtmhMdHzazLMvkwcrx7kTgehUeIcQcTWowrf9yZ1VubmfmN1N
aCorB1S4bUHBCl73dQgaKHm1HvxugLb6U3a6SA3Vmw3CtkDeWXChid3no42zyM2M
XbjOcfzMHjqCBCzFescRRMgk21XXj4f5QUqLes6qlcUllxvuvpvfwpmUqGc0h1pG
fruho9jFWa11ensS0DeOUv7Q988avnb3PlI/gx6cOSPskiMki6uz90PfHt5mB2za
D3vfpDi3qi9Ixrxou8aEOcKiPMgJheekAfG98pCwsVqEojWiZ2ijHGKy/dDgGpYx
KT/3FvsmfNOhSeuVZ5TjwohtFEyf+APOKqfbvMNOo8ILxJTRuuRk+nHqoMVVW2qE
jFRjuE9Hju0FUGiZcaJpmKP7yTd3hw38DkEsbCNeg3WpnEhsWzXW4zq+ziacrloR
C8rdqmbzsdx4cJvKFU6auensnPurcbjNImlnmKGjqWP8a40AgH8K5izkeYr0J+no
u2ARmgf+5+N5hRz11XsGveUHLpsSNnConbM9aTc+DakOQbOexAvLvFlwlrm5pbKc
n66LscdHU85V8RfFj/GMeybFXe4/5aE3jkGkxUDWP/Rr9inlJiZ8v8puLtwBiAk5
+jYZdmpbYs/YUhZMf3cND0Fvo66/POUjhTyoWgI7yWrMlWGFJl3fp06iNT8v3kZD
wuUw2p2BOY2SiYv0uqqZx0Un4B7xZQTDA9GCVc53fr74hFmzwXMqlzP8nWSrQ4g2
jjnYZ4mvLLP8rDgbw6+x454ThM/5mdCvrnssGIowuYmdzn7uoO13QL9qOE+KD6NU
2SvbQaZmaroPFOCFikNHaCHF0sz0QxW0Aq23kqqUKp3Sn9OGPpsXtjblgv6Z2sqv
RVl6sGmzSqsQbtSFn3DfYOrqsFTtmTDIQ2+nNdxlTrXJAEjPZS8EzbZTvggdZa33
kgGBaDe2yJvUfowiTAry2NWk5b1Usd7xuokmAGNjizxsE0rHg/LJgzWM5a5rrEaE
FiVCVyBgIsiUaHPRkvmnEcCQfQQ4KwTm8Cq00YgYceQhtUryJ+chYPsIyRCI0qPB
wWbUBWGqHPQ8Nz56q9nKz/AYc3IvaZXhHDVulfCL9FzBkqWEhKXllpUIrx1iUj2d
WYhLGE/umz9TTAaKjdOA+OSUw6SoAbcXv/r0UXdQcnQ2sDdq8C03Dc1Lq0p3n3Gd
Eyyo85AFPsYj6LzzIHE0fNWCpIM8pk2ohWJ6r8dKO9HWusMDdIR2/ujk8CnNoyIy
Vwp0bkGnm0w3tbxwEqa1ysN24waLO4Q3CRFAcNyl/ifMRq8IKXnpzM4xf0TSJxMi
+YFYmpzRhQ3lhtqrRJ0BtIDKuGV6auH32YVX20JUoD22Z8ANg5VO7CttLLrdalgO
TUbGqIiRQReofOMp9OJrnsO6/BrXI6KKGbwREKl15kT9tbREkWyHUQbYgBw3U5j2
B/Z5F6c3PW9CSyW+Gh5y7f4S27gplI9tpsZKUQMK/fdwFDq8JstAnvVN7rA8EtJs
sTfaK8pIPpUy2a+AhKGQ51DSGYlDE1ld6KPvO93wgAEMs6phOEyAL9lKMW+mvbGk
dc+6Eu3yWgxbNXxgVTJYVz/KaBL5tj/wSfO2CwSAbh/eOQMG9GJWKsFBHpxom72v
U9T/qDKujFTpWngyO35wMCTozE61lqaZdhTKcLQmwn5cu3rNdVrfov7qS5/foeSn
ZVRC6sKm4d++KYQibnr7e6yNsrxUJVVulN9rSgkpV/Hzy6v4kaF7PtuIV5Pb0eWi
H0I6Z+FnpwzNpyOsDQw/LUzMriPyAGigyfMv4xEpzA9okMdk838cec5vIPS7muSM
Xjzk7xKyIFebgEnf/w7WO7e+E59hfSKqsESP644/nd3A6KOmf41rXv6cU5p5UT8i
uu8/SGUi/w20uDS6UXwCoPu+KFo5HNj5frngB+FwjXOmyYLTAeMoLWb94fqs88R2
6uPD8kS3itiJltJ+BDccru0eedYU52oDlhpI/zhYE5BXh/MQ6JZh76uOy6UrAfpZ
pR23slLCcvNuR9AkYhHhwlbn06wH08nArA4SPqzcZh60mn/qzD2B5cTdr1iJef5h
kdYRAMj94bvIXPyAJ9a1mztdnfT2+8n9sGWD81YkEMu7P0bRLpouM08zkUT4sbrw
2Zvz/swlWsmzhuhrPhcOYfhaeIW/+hc3nhtRUYPxec0YLjKopKVgwHvtXMuFeez/
qkBVd+4WImm4K60Zci5L5PPYEZRHfAIYc+TPGQPpvU74PRk68+Y6bkj0byo9LIuV
NRWGFFnnHpdscp+cnVSUCC4PIb4V59KIj68kkhPKt0jWFaglOMTrsg2WpdIZDDR4
UcuOd0mh2e1een4LJNLHodBFO+eKGW3nRgoqxBko2hiUf72qjAnq8jUey4rtwsLt
QUgoypjNnkLG9ZFw/0Xga2vKKF85GACS09rBtpsWczuA7YxtqqMwEvcLQTNNYvrf
xNOoKuyDPBtdnv2IDu//pkbaF00n1FynnfLLXO32xDbvPgytqME4qww4qXpL/vdK
m4lLI6gty4VoWOlxr40GUS3yURV6FIosY7vMF3z0MMrtN/5IeVtX6WP1G+cdQGJv
gH9bB5J81hTYrp5bGeByNYLc7bcbf8C+bL1EIe2EqqucucJmQdxsXPN8rPMZKFEC
3M+STlvzOVw3213la55g6bRN4XDVlW6nzta3ejo1o7+djfAcuvaWAag2+uXlc2+3
uuFguBX0KZ5UWRj1LHhF8fiEnSvg9/95rZ/sb7236zLpoj9K3xxM/AMB9PJOi0P0
zHh/7Sr9V1yD9ob5CU1gF1j24C5cvu5Mo8KbdMhxbIOQXN7wMPsAZq0Hd+3AcKbB
/AHEGoAARD7EBCw6i5l0z6Ou03c+egakt2XP2Bufwh4bPC9NAknulX5alu3xpkFc
W+mk7VRjTEXUKKCh6HtMcNT7XR8bD/+V0fTQvBjmPGlTr1XlgNLm8bl5VUKrDvwp
ZK51BJRThXGNXY8djlSWtHzYdBqQd304DSs+A9A4KMVhFpsXB0tld2v23QNqvJ3J
SqJ2wCf9m2dFV5GIUb+5fZi7HNtj1Vd6jlKJvqkRIB1fpfPmIlrTdmWfuPqVpFOa
+2kNf26NCXl8sb9euI3fB5oBKzQAdeEILMmfgCPMMs0Rp9PkUu9CFHiEdqLwpaA4
ae5TbKQ36YQh3IMFDPYkeEnxYazuTovJuSlDVPyuR6tbO0TATh+qZLI4tu69oYS5
UT3mwzA8oXYCsCVl4y8jF+MjF9uQcrUOlo4yek4a1NVh1x4E3vGP/v41c5RBCeYD
HDeyQ6T3D6xxW5u9rSPR+SVs9fhkTklZD+jKIzzsfZSgpupMf4VRcdltvmJbuJ4T
OcSPM8BM4gZJtAgcwbztlGL9872EGAM1ILPy3H4pKq0pAG+MklAvB2HjdOkx2Ic1
7GrZ58B3CN1oRKnt4gfraa98yFqG4pPCjCwAKsF99YJf36HCQ//aVQyby0pVQOu+
/qtmTpMRCa9KQ2ViHBqdzLajTAthG88Pug47EO/86ubBj+jzNLqGYPXqB25BFLRX
PlhXlD+uXiAWhhghS5ZdO3BnmJjpehXrP9NDD8CPc/VvPXUS8MaKSrnZ28NE/XVv
HYMjA1KYq9AAoEEhLx+4lIUtm77z3jkS4Xlo4oFFZ+mcNRrUI8pgfsl0J83aDk9M
+AY4SONGEUc8ZwoZ+pxjY9r0xrYEN3EgQlXdyKDCyAeV5jAFeRS2fUnCZwHQz1a0
3+tMIAF6BpD1BHkx+uP+4OVf0zhq14yuH+bhYEKp4CiAoiRFAJc6geVC8UIlUg0z
BpF18ffaLE9mmr0o5sQr8Gyo29AdBKIb06TBSTvgXXaF1bzt2YnJmSI5fUnvu6wM
j4bwebGZMdgoARDBYsgAOx26uHoYxmGhHBtdhAQ8YanYy6ddkmkT0cJghnM3KgxG
CEo9U6jOzMvSvbZbkbWU84BHLKoVzm2Pi4UFp8yK6kQdg8jp4q40+PrPNKny8qIV
QLDwlWSZyL8za7jGMOhtcbC/QZV0L4xRNAjA5x0eyo7Y32sWVFmNuOlR9YyYwg+7
cpUdbaC39trn1AaLEhL9zZlzqnqjR206q5I5+YlOZfWmHiBwFIWz0/GklhYJ5cGV
XOQZxLCgfN+d18hbIrvhwy+4R5I/4AfnOGheyNJD4zWmBN9mZPDyEm9dEJb2od0R
fohOnXEFxPO+W0k/bNzagrgINNZLb7MQnXxUVPjI/GGpvqfAXoZecLt8D6OyNagw
nO3mhJMEsfTYzVGA8rq36/Za68BRmZ/6+yKKaXHNfgjmOKW0FxRjK+M0L5sP+w7g
Gvi7r2H3rDHjzeyCC3e5WLvcZTq6IZawiRJ7eHXw4Th3AeexTnob1XHrXZ+XoDRX
fvjWjNz82yRY7RUJ5eau9WNtdHAeeELWqBf/Knd6h2Ci3UTJLY+gd0xc03BWz8EI
fCzh2C4FmLC3VahIS/x3Q4rNIOVMqWEDKpt+oZuQeqYSWHfUDaZv6TQtoV/ZCi56
LydyiKRHLYha5/Y+xTmSYCvnmAFbS/HSLNifk+chPqIuACvT65+V6LvP5X63Uk3E
x8ZbYyjVeSVlU+ffI7Kt+3Ajs1g8MFXhyKLjKqxFCuKPjHHW/O6wkkF64wdwsjvt
w1w2MXx9HYyd3mz7g39/BBqwSLwIwrEELbf/UIpw2gEhas5sBm7C3KDj/jlKrEL+
wELt3SwZfNLV6/ATXElJ/f8/a6vGmaZUkADc+S4VKcXRsgwKf5OFhSYg7+3IPmRN
hBClOSF+vfx2Sg3+oX5+eTJ6oo+dkB6yGzuKBDf7k8e+OD7woRL1+gQ8+nqUd0HJ
a7GaFraSeB/Sjj0Lqmz93SJ5z0AC7hVpcxOOLpwzoJwgAmq8unuOB7S64bH0Xbox
Zza1XNSi4bNCj5mND3A8W/TSQwWIBd2thvQgygXSWYAsgsu1ih+rupvZ2x/5ul8u
/9VwqBp6isnHe+UwldmNBz4PwDYCbfxyZJrDZ3FkDf/z6xSHg4WRB+7djk+cDiCp
6cgpuuU4ygcCLSewHhhUbkzQfO6Jtj7rMLPOCvibkUxJcROgrkcoZsqlw0VrTd8e
YN1DkfFfrbbxfvJ30kXve6UIeHBTD3BXPzxRrU6MIpVuJPK0B5SWyADL9ZSRiNw3
dInx2CkNLxPAPYJVqvBx4WvX+2ZkYeli7KSyc2nHSkeRJXw9WOy+jKQqiR+/MKUm
WcqFIShFMiU4cr4eJHMfbO2vEuhNtFSOTng+uhKobtGV9mQ3ovJeeOtHJXk8k0sl
RImZbYW+17FpzsoG19Go+kFWh0ZS+fZ4oVZXitJ4JDQ43dbXKm/oiQlGEeVKahTE
sDsGNMU1SxNv5gA+YABvhFNxe6ZT6uLxIb4W2tfL3KDaYg7QSTpTjyzZ78d19km8
qzCRIe2amHZGbW6FYSJRnXOJzj3dLRH1aal1Mp0KJC1bDDoBAsyvnLLe5bxRRF+W
q3OQ0ZXmrrvn7dYwJ+vB8VUhNyeNKYGiAjafi+PUK+vhyvKTbbK5KciTc8UQ+cWw
iMB9wx8BlweIku/n8XkRtc9PXIWbsEnO7OPT4EUOnzcB+eq2mXVV7vGk/G5p2pQS
LyV8vf/7s5/7l4ULXCQqhOcwulV+syj5+RT+tRHMn8lP6RDC9ypblVsDsv46Oltp
6YUb65aAn0kP2WQqzty8KDMs1d2/M/I9B9dB+tHKnBxrs1RkWh7D4O+9SoxINV2M
CzIJNQCC5IhJDlRCA3e16A5G17xpYowzuxy1dYq42YrYWgCrdtnCfWLa49QMG5fz
k80D/Ws/6bQEHjWcvncDgROyoxTeKNCDrX+5xaMq4/nkbUxrWQUDRHfQAZwERY1g
y5WMcYZSfZ1XVz6M0ZXPz/8TPdlQSXSRygbXiiAkEY35p4TwTW/A6zPd87FpXHe/
nsRazp4zBvuuJ00i57Mo5xUw1EOmlSpZq90aZ/0izFDSZcVuHp1xQ7NOn95rHAfj
UbSvX7WG/wn6q8zS1xsX9RQlrLLwiWHWcafPfM4Qzc69ugxSLp002L8P5UsSs2js
17FHSJWo3PXdX79BRlklB9F0WRl/NbLEas3K5qOpEy5N1646PFi8IX9aNiHoW0Z2
bEBo+9BJ7e2f1/kz6MKvJNl3RAmfTxxELlVo18ZzXgLICfpj2SWFRqp4JXLhRusY
uFSBVwT1GuoY2gGSR+2QUgj/fipXSVt//MbvgyuErYB3nBfAFIxPafCa+JBemPtX
QoZ8SO2AwVIwhFQP0NfymtsBfBpSak9vJXO4hl3D+FeuFFKMAc5Y/l2Odif0G5BY
4HJUStpNYFXGaJSOPnvPLkA8u5g3Szq1HjsTBXyIFB/IHZjZSX6pOgdXNOcrUfWb
cuanJa6yCrX1EJuwAkGZqYInVViy6x4+IsPhnVhRIIptAyOPaR1lyeSPpwMW5Mjz
bYk1X0T5lWaaV07BGODZrlO0fnWWGxRBRqO0NrWfD0G8plr7G9UZZEgDeXuPAMQW
rGJOVHyYT8mM3deGsGvbpOLUafYQEoc0tO95QjtazIcDG0qC5ZA0eOXfAV7o+ZUs
MjtW03jNllVGOOfuuHZEHEy28X+ksNsJ7zC98OqUdPw61bH8sl8pSJVBb1DEFZls
ondmi5C9aA9lHzq0k/P194MFxqETW8+/SSCqb4Xnn5J+5C2uq1QlpnJY0b1eGclu
xyKRn8yj4z7h7is7GyDjoV0mnsyq0L7h1QLdXceYcHUpl9Thz2lCYpbktm+kVMus
X3JG4aV+02CBJGTtsDScCxzjuD8gBZ1kw2Cb2k/qG+9OLJiuQ0FN4yvl5RUrJBsl
ONdv9bonTgtbQ8PnZoIrzcOR+WKpOcL5fNU3xXYZnD9UKtVrkg/lJeyAIuEVP6x2
uQfepaQ4gQlYoXNOLB+zkYMUv6sSrFIUUEcjH7D/6bGg4pue2Rtw0+Q9k6Z8FgEp
TdldPwBAY2RDU3q9c5z6LffuIlyBJUjtFbhTo44fKq4Dnwl8iUoGunj7HWTviduP
zMcGOE6YrjFESoXMzXn1wgzgK7XcJLYzOuM9gBK2ssCk9GGclps+g7b1Tse56R7I
UKHk0WocBt0EubQERtiyDTuknl8INnJSfREJmdClEFoHse+KDRlZchsEimokQvPw
q/QbK9DmHKWrA54eYTK+01TJJ/FfOahYDzIfV3YtDx+lEmqiwYai5Re/EZo+R5eo
dszijjAIWh+qRLPhgiLwqRxJ9JTkayHHor8JTMj6dy+2C1lDFIVMYGyUr52Cjvsc
Bk4Po7oWWpyAOgOWueQMLgnqvPq/6KEqWJnbTjjigT4RF8l8LLdk+zUITUqaXKJL
5hsHPAEg8y6ypd+QOlm6kBRrKkUTMlkhKWFDSUX9I3qkLZcTMRhfL+9OBOPt/3Ye
IYTX9wcIA7dlawT+00CESCx7rFf10aXuAcbxsTo4ukgdv/eZ+h15yH1gdvfQfaW+
LSVsRhtoaSErzh4j8z28qcA0OQQYAk4zJYuSw3EnUOPVWq2BH3BOi4Mu+5C3TBNy
askGwgTgyhnWUOQl6M7O/hJ0KArqM28cj7lVOf7vYCLtOOpWNwiyyzFVacs/hsZa
YaPptw4EQPJToicu/kL2+pzvbekh5Ds20Tg8LfGvZw3lAnOm2Ft0j40tZX9IzIix
W7Ja/ZvOb3DsSOitWes8xoFlmxyVz8ZSyuzSpU2IbKJfo53I7BL7+3w+1hsmToHI
ndSFo2aDdtj51Q22cKDbVc2xdDm8MziG2J5jIio5Y09P0/g7h/ljtzIMk86WCrUD
KtX9GUe1J1l/7c1q7d+msW51pT4h3guagcP2fm0Q8kFHciFXG5pDYsSJXKCDpgtE
jE36VxqyTgm9vtuo82S6lGEwd8g9MHVFaS0N5LXUrsCv8KemuFvetWcR5qnhxC+Y
brz6jANJeE4BWh5w4ui5j3NKifIuMT2b44Og4WwQuzCWdWYf6XJVuGttybIX4vmI
4Oz3JQbQiKxQb3X/cIMrxYrmHseviyIX+I1J/Ao/rXNVt0/xQbyU6r+/QTVD2bMK
qgDMvP48S9J3peqnCTWG+A1eKfHPPQ9gLGW7DVi+DtSakENoOH+kd1TWlPXn8fnn
h0k1YA/vJT3Op9AFe3jPXSyHHTtKVyY/eiy87dXmoFfI35avw72jFw4peykA9grj
J7zescT/I/zW1KEAZIaO0+CKTtLYXjse2BvvozgfLHTN0rbsIYLVmH4PRSwmvx83
rCJ11KuNFE0mesUfm731mB1iJ6lRfkfTBG5No9L8tvlwNDkqWW6Jhc4uH5fv1qUt
NZ6vlR0VqK2ShUEHoOCZapeD+x4ZsxBHF+uh6Lmwj+uZ6zyxJREhZro2auNeWWYi
vXPrHd5+9smo1DcIqfqsMML6Gjk+SMRlq/vVPHZaIOJ+Zn0qPyNwActHquhiN0HV
2QsjcITPFcB4mmfxfb+SKmiLs7rmK25cHyvL+bu4Fx+VcHiKpoLW+CaX/gxkda5Z
6zSgyrlagTGV+5oaAIrknwvgSAnyMg5/uEWhdksmvquWiTECUbfGsAMdPd0nD1Ej
3mt6p9PEkWrUONyrzAa8DDgET5sczxlGguNgyx0KbONWGB+zsnmUhC+VeEDWSHhC
Haf+FLVHLpuqGwoFqJH3UnGT/W9cAL9ZI6JK2t2otP4+L34m05/iSCWF84wGqtwC
v42HREL8y8Z+nT/Q6gFkToUmpQ0JWk54LjnKSO1vLh08N8aodwCDJgRjNEQgFyP0
Rtg0h/pUopSShHvBSkq94mP2RgGz+N3g3bDv0RFiDlxt91/wO4S34PsxlaIqpY2y
T4uw+W5YHfKxStIMRWyRKtxuzmYKcywmTcVDTdxgejQYPWBoGg23njODhgVoScs6
ray+7J/LAMM+bZjV7h/Tdt64RJT2ALXDKTVdNoDjwp0whKpf/BK0y1UvPI8Qn9wT
e71nrhSsBSL3GPxh7rZ0E5IFsnadNB3E+tpA9ow1Qb5tl0tltCXjBs5JANq46JSw
tbY6vTKzA6Cpzx0d+Cw0D84VukejBMjdQT5fNE11VceT45zR55lKgjxsJRUoU+64
kVnk6VCHT8E3xWQoNlBjfIwVnpw7MTu43mA/ETkLblkfxtrsRPx8BXt7pCU+DFYa
iShn3R2hOQjMPcVUxAU9RcZMoMIfvtIOKjZg+OAspnlW9uMupxk5wOyUeGeHk2Kc
mGJftqOGp64sFTCcbz/pxyMPwDu1ocy55y0Mpz5Jpo3CaTP5RmIu14t4aBUS1mNa
NpKu0+5HsIdKvuu/Bh8RtkLaYPqzX0rYS3wzP26z+KFHxWmgCbsE7bUXMj56/avo
X0ubxGPZPaZHLLFeSBOILCofFqFXc+qb2nkiycTPk10M3YDN3G/cxROgnfW967hB
mMgMbLdLYWc9EiPo7N5zD7ePZZ69PV3I2HKnTuW7i4ofszsuB/sGqIVVa8dbDghz
bbWSHXn6eYDDomih8qMVwLWnMQMFhsAfZ+qxnvtB+1FQ7jKEVt490tgtiZLyJzlX
4NA4BUSQuxdAU74KYhvtMoUfc3SrGuzrhr5rN4fE/hDGwRG+F+lT3dvioWxqvx0s
OaThaWS6rJNloVNFGfIbvzjMLg8TZRLaFan/Mgf82ohUNrUurI3U7u/algxwqXdX
vxYjtbYvUD8MnKOCzpV75QlWd6Zz4HAd48kcL/LHi9IHPbr1mfpR0AfMaKaq04We
UVyJdxzAyCCuIh3ex+Cl+OCECOQxTtjv5zwCDPyeEAjNfliNFNvZD/h5S1iCi1KJ
eaCUuNm1R1nTUBp7BqNYRXe+pq7xyzkrQc2VsFVbiVVzIVeJpGiDMj37KKIsDsIL
/kSB+bbruj8U0MxJ5NkQSU8I0/v4fqlkYB0rs9wVpgSqs2iRHlHM2xyCZ0X/dVmx
YxbpBy9B+Lx23xx3cYntiX7QdK8NpGqcKk5bb4GXozurVMv22OCCOitPrDwUizXK
1BBmmI/Whj9sJLm5i27xvAt4gAIBbkuJEy4lYCnizjemnLk4mbQt/+WP9qTnwkOd
yvokfqngAWp/YpZ9ylXIn/giKVUiD6rMcxsGNKNjTkI7gNUDohSneQ33iVqBy/cL
KVg9aZUw9vEaNtisLaYec8ms5UqJJ0o/wMuGBsKi8eflueJC9J4cy9y+AKYwsNXf
iZNUGu+KrCMbNIqGxHIhSxP37qKQIaN1wD6oLgxhoH2elLpHZTOYTH4jSbp5R7Zk
pEEkGJWixezZax0d5LJuaKqurw85y12BX3HqzjXWpfs/556vC0cPxZhozQS7p0e8
IbhGbkkJQLUbMZzkNf/OIPNqdaHAKLKy4bT8UPO5zUHwWwu5JLNdbc+O2uSdweOa
cnDbhtjoO1lEQk0eQZ1v1TYh84hoJ9pD5A8c2ZaDVFdQWxme9k2UkhPL8J5cjiBE
p9mkUcR4wKjBTlMBX3PwlTP8kN/GYwkrwubqPaIJCqRlcC32koyAzp0T1oeSky5a
zHpZaLiRv/peNtN1V7RSrSqp5BjFOVbkDMLEe1eqY9LsfhixEPsj6VL4B2Trlk9q
6ZSDKSJFCZLP/kXYS9/VCDJ2DezOzBr1J1qXFvdIE71t9M1jgD+PWYSB5m1UUVp+
zYgnG45gcrHIIuoelLN+vzEfiFtCyXcxSETsaVFyYX/UOGD13BMiBl0KHoghnOSm
8qf3leO7f7CDdK/Q1G4YyVSTeIPsXsL5JNubWDaD/ebbwxcbsBuybcLUQsHz2or2
OzkSgcm8y13V/q2PNBuY1cTTT3jA7/4yMzT7vvrPTirluqH2x5+V5Vus6Cc3D7kI
aL1aTmMNlinwBrmd7fI2wu5SRB0SWy35rve8AZMHPjxmVORxUeTRQtn6Uwb2ylG3
vv6ucTvCcMatPkHJOPWYbXQRq5nMHae2y4QSDLc1Nj+Qu4doxrTlQ7ynhNIDJeQk
PtTFk4YBED0FPhkrKdU9a4dtm9bW3BE9pykCPYIUGTEnmxQHpn1/BOnzvsjm4c9T
BOAD4OSOXahcKbAoVtqhDMQrOy2zNfCvM5yXyzOVqauDh9fhrYntMJdfrh3TrWE2
ZuYFIu+iWJFx0tuZSJq5F5fpBC65N67xkenj/4lqCQPnsv3vdBizT8sSZQdPDX93
fRTpsarWIcLnSpsvjaxtC6+kG4FMPpB/+/4ELwvjLFQaBWB8ajwJv29zSp0yMLfq
no2R8HUfayo13BNotqtW9Dhl5Xn3pJ+3WxmPUzlrzxqbHfCiuvb9d3NZUoJ/CoXB
L/SLZBjsSkJ2pejIiKfD9tDcdT7RrvczHkqnob0E5cCCLMVIfqDqAepYJJPQIH+i
F24MDPxXWuMNhI0Z16/+uAVwlCIv+aIPxuzEWSp8uvfIINavHoKwdKIvD3t0+hht
19x/SnDj/2Ak5VBrfgFUzQf6mMPEbsyHovx5yE+AfqP7kHQFMGdIZ57VxWoAwU3S
IJXi0YgrF8gXKuaiYq9WpHKqEf4/GzcYtQfEO15iGw/hyv7s3JxkZo5qaX5IKfxx
HTgeOCxEdRYv3oGYMq+B42k6rgKy8Z0kytpLQ7xLIZ26/KeTBhjkvVIg9wC0u6ET
3+3uskunKqlryCZTTjEeCfYR5mhApSOCDM3upfizDCPe7aS/hMMCE+aXXH4Fg4cz
ww9dRadHhUx4+9KS9Rb4Ug7eay0eY1c5KkN+MbBavSYR8qZ5EFpOKsST1EyExl7O
yHdqqqaP0muk5Si2MoHdZxQ6pp3DZ9hCH2rtZ77YDXr85t6GHZ203i5uDgoJhrHi
aEFvFAee91mdnxGIpTes9rAwVxQU/rPbdih7PrV9LmcqYbevohdaAgEzY0eKF9Rr
YvIH/0fQgUWpkylg/KMvoy87BeXuLTbE+ZH1gE0XMwaxGcTTfQfMy73e8nnVN6mC
GKvJjUyqV+PKNkTFwshWEOjVo86taKJvjujND5/3Oqi0DSuR/Jy0C7AOo+jXzFGU
iOXWr7E0las9Cjj98/dmbKcyP86ZEeV716Cpolj9rsobYpyT8igWI7rjR+lcpIvu
fDXFpQM3cdoKTIKG8pBgKmP61bMAqNqU8qU9YCKona3umUtw3JXD4ScdeRShslyN
Z1M4+mD4Ir2RvuRSKoXUZKG7ux0GoAYgTVxQUQd1/Qnz+J+yfXJ51dxiYwwuJn2e
QtjbG5TIeeOg1sRzymizsbEaBse2MrUgpYN4Nwxlg6ltsaCbdDjg2uFplKv5a0ab
C0qE33gLeRsn5tpVxe+abJ7VxMAiFLCbcymYVm4hyaeGZcK6HU+9td7yAsdCG1VW
vkKRPw8mqVCjMw4yefnDxjHgPQB9xq1cHug/WnQbA911yHS7GFzXn9WQpnODSJXs
3O8sn7nzUnopRxo2LtbJViKstxnHbTAr4Z+biUKSsurvLpM6VipxBPsnsbHOkAOc
p2Rs1y5whzU/Fu5dy4xOBgdmM1iH7HT/TYK5FMDanq8k4IM4WtKSsNYCnuHlLpw3
rDELFouq2EeD3l0zhNdyFHVtS8ZzZe7u59unSksNgLKu/TTUBrp6oHgcRfUm/0nO
iftyqHQ/CRSmxUR4dlzbACBS0UMhjmIQSoPTpnwahUEfbRbVYf0AWmprXIdeohPp
sF1XBJYEBiiNs8093qpZzfojnrpgA3cBSGarWXKp/i2R9H+/gWbHPWposjZrB4hS
v6Pl/R8g7qFkrr4RBpPPdvAm3IcxjdCIovRyaEKKxviDNSrHog/xiqb93EYUV88t
ovTJpSZYzdJ3HUC7eJnu5vE8+34HQoDEdN0nirtLBYZSvK5xCZPw6YEbMEul1FAW
aJ2iUcuKeOCX5hF91tpRc/ZmOb1DpR6dIUOPfLtfs0n+cqmH3W3SHLBOTWCcpoCU
yEm1uieTx8bBmp0cFCIx4w9cC70Y49l+4bxoiqBsm8O76rl5CES3HCwPCWwL33SS
gbMLFF/SZXFj1/3/EfIc3u8QAB6hThZfNVt6J6U9U1icKqmnbrPHZ67gmGa98v7d
HFR7HEmMceFvfI+rC/4lZeyAC5bNtbwmyA6XF50q9Dt87bb1PcBryWBI1lPvQw27
h8vdgUPA+WCFsgIXU1qqBmaSQ+ik+QWJQiSZQ9SLQCHMMisTjGrzKeHcp1lfVwCM
fw1Mwlz3y0rHvS1N0aNisFjTL9h4o+Hxmv0QEbFmh1H2/hDeXEPc8JmZdh69WAOX
TWOS2ELzirxMRMJueFz7mxc8hnNBkDpx78d9l2BJBUBF2Z0pQVv8i0IsSEYeBvdz
dzJI67302qaTGZtaE8IatZtMz6H01tbPhcmUZlIPCHWZfvKACRx+4TEP8nrcXRLO
ekqpY4sqW8dNX6w4q8dylGfstIEnYji8D8yvGS1/g+RQSNR6+EvDUt/FUDz9RRgy
lENVc2JA6YX96IcZXZ8TO5ijPShoNsUR6Cb8t4GYbQA509HylPMeevA6WIzj6YjT
zhDrwKdExmVBOocmChEkJGfeSGB+aa51M1Q9TomQo9+7AIpvq75cfOGScITsj0gg
dd9E3rMVeiT1VT/lm+PFWlZFEPTWhjgEJhnY8VHr0HAo/EM+nmhqgrQ/wBVZEN+U
VCnQzT8sGRwfmRFTsfXQ37a8rftb3jJmcPRyn64B9gAryc1j0SdNOgmuZhD+8My8
kVqtNZRuZEMCLCNdnYhqm7XcUhW1unZl/YA+hW8AYJUxoyx+/epK/4py7D+Rs+hO
SKlvcf9CG99IR1qsEd4kVaSybnj5/bNRpt+XPna2q4E4Z4igWaSehUGDQlBVFk0C
9lr8+Wnrj/jkkk7LPWCewqQGeB+NUkmPKF0tb510ZC5en1Jp/bnxSHaQBcn/wPSP
+8v7SZMjXVnbBD4j8XHRn3fHjaJ1koZc8MuAgHJ4N7oRIDTNmUEE4JwcxQYaWAbu
ch2RjeaixIrhiL2m4nwzMO2We6qvZcLzhV6TGFqTE5rvB9xJeonIugyN7zM+o8AB
FQldkAeh9877FIOClUxsbxepHoMWnOePxth1dZ79Z+5cIkCDyJdq849ptxcVFg7n
kCysLlVM0+1CcEqy9XitDib+1XQ+NB0uY+QB6u3hDuE5b8WUOq0kQ62vnF9tnVGk
sl12c2zMqHlezWJqRSJwvmh8WmzVMKH4e9whCXSgtr05NliJR6pfSfCC7XK8M1bt
XnQtvTi2ZO3w38O+0RHduhEzni0LaGaBLyu5HcAkd7zC3ri2Tevyd1yrtACMJm1p
wStIdJsK2REfdxeLjxe4MbqCRWA6FcMS2vTA+OhbTm9gkTl8VzlboothPPxgbXn8
hH3IHKk4F4Ptpr05iBzlUgB5kXX3V+EcNKK1oYuz5C3nfCBua3Wvs16hzPi3ESAN
t6a1nFTeDNZRN3WMWXSa6+pS6anzhC36jDQQFBIAmyRn6mGUlaR9dEZDwznFWQVL
RMikp4GKtd4PxSiiwxAKZeUcWAqfo17jcAphFluYUnAEK24C/35/7cj0HCYtPan0
gxhd1axKjsER0cvJ+eMue++YPVF/QMkt5/K88Lafs2zteseiLktVutKGiI1QbMcx
Etmi9/Be/YmcoZYIJ8ywzrewKPXTMbXAhrHOmguMkGmWWcXdbdrQkAIwmPqg9zuo
EAFfNc82YbyTkDNL54ouJ18kq/eWfSafeQBwFpu2N1E+kMpdXjJ8/HUThPkpRZ0W
qYLyo/OiV56//eOKoke8YrO+Eq3e2WPavQ/Cf+MF5v7m53J2MeGIG2Qf5hdghgJz
QUhb1IlRXcAWkrnP+uTq0PVFLIBGB3j0VDL3KaU7daT1NFBbccCCqYQT3nQxu62G
g1JDMlxov5jFDVSTX8SBNmqgDplWjRckMWieBS1IB8ScrHuI9S/7/FSz+1WyxUUG
s1vIpmF+OgA5KLP50VSej7b1/P3NEg8AtVYuDrEdjCNwLYQ66Vd9YYE6TGgUMZhJ
vPPoliadmLQj46/QBpIpG9itskAazPBuaIVPFd58u3U7V5k7AMZgdRGxTTOeF8k0
fKCEL/ZviXZkqFL6GbkoOwjWnQZWRSdAnECRBHHT9gIk35WUUbPfKF+zB4+VGIN0
ue1PTgGWVpJ1Qz+NV4kpny/hEq4Hw31exKjKK6VkVLg8JJvQM9iMbfI8ahr9rXU9
uKAcIjKmGu7oSO+uvM40YFqCRWr/FDAmwYPShaAGjA9MdfEAwe6+zfc4cFP9INVt
sxTIoR3r7aJDTvvNt15XZV7ECflPCs2j6z7HyUkBV3UA92Kl6qpif9IG7UOGFUJA
Qy8LFnFcJ9zHcb1J/fOqsVv+ivGNhTXSoFKrwzU8S3SJUM/U7GGMspgqO4EjuRpG
tf0Vwiyvhc+QA1V3lp98SEpMkxL51Ou5QgVaY4LKn3dCT7dIM035EVF1K/tYxBOj
KlJbMeC9IavqtF38KDNADRmIg3iSPIjWuYFCKC8cQS5Kb+qaW6ZpVGjOo26KGM7N
IrjX81rONuoCdUPPhkgclV+tHY4EwXTGt7LZ8HHdIclx/rONUMr8bCfRyXiFloEu
WgGoYbhS+YYEnBjK9DZl0lajyu5/NPwXj2pFNDMkJ1GSmBglukYPvQb6SioaheyW
XRkmylOff0P11OgutVCIH8I90HfAcMBsFli52we8xvWMWRvmagze3xd8AF/4k3lb
MNlneruPXuzbnJOAxCDkYvDRCxtgzNfXQOXyO50piCazyNU10VOkeEU7szhnwjpA
79tBvJbr2KmbER23eiXcTorTILo1BFxD3RuC+OMl9lT34IfJ5Qu3zw1ZpRK+jdz9
miNj3GJ1jY2TX5BGwat1eCcJ38+tQB/rYXCHG9vcL4SkL2TvRAfuVN7Elt98nKjI
dipS4EReDLxclfQnhIdSQrrVethACL+H1uY+DaWVCGx4ZE2rnYXSr0kCzrFOy/u5
X5kcbcl0ApvVt7gUKwqbhIZ1lcQ2QkIIvxvNN8ER1MYZfDMPWjKeNY01MfLzdE73
ZTk520e14FJtVwLNC+3Vxc+BAj2U/W2FRvbNAEMhI6phoNWN/EeeIn2TH1bwDr/y
9YaWr1VIiUTZ6P+7ZJ/DtdnPychh4IUxNOUnyQeHXn1341df+rgOSHeGr2BTzL5i
9Y4bis/6f6RheUhYYB//+FAYRqNDGImxNG9nZHVf7b7X12aIJFea0Ty9RkVPLHqg
Icga0ZKXQRP7mdCklhFr6rlhZ+UYVyq2iJYCcVqXIbwBnD/PbmE5NJ3arUu1SXpH
HJAHkES8SUoRXIXFyaH2JO3ETOWsvvWwuWoxEFzZP7mM3+5U+eqJzt1+YszccrOn
KPz2xcR81eoScTJSOt818jHDwJS9p/h6FC3BCS2uJcH7hUB/VHf3YU+8hxSHMos5
IDnFU+GkSsaTCUYnjy2GrHcnvrxZQzg1pFugu8qmBZx55FcGHKEXdIBzyA1Zh7AN
eOJw4cLCkB/2YfbfDnY4wJ4REg8IYD47A7F3poJ1af3/zIZophA+fA9GSeIJ+9nP
VuhkjyQgoc04XU4SL1ttJHXHPBQ2HRviPPH7eRB6qy9MSRoca0K9FHMzrP+ztgvt
cQFRcc/9m+rS3S0lsp/XP4tFt03wVaOFi5PraEOaH/mt7eGjWszLvx0wpZpkWcSz
D0d/KEmT0QlF3ty0jrYhdINdI/cR9hWNvGUIQiZTdyEb0pOAj7enxBd6T8DQVH0r
TI69YZd034wEWGKm+5eoTqeHTCoH5fGbKBNqExUJXmz0LiG9Is7R1QI9fFOe7tOn
xPMbl/o91ETCIjdwGH2EFIdtwucKNQP/ftcIc1bhKM33x8HuZ4WmjF8oNlZsiSFJ
EW8TZGuJtG20XgMuuqtaUOxq+BR6IYn1DRG/XjpbxW22uHGqe7p0Fuu/aJLGMYck
u/heYYEQ5lSHwEbkTrSvKaygqP8yNEWkbziZUa1UFe6YEqTtG5YlPxaqGzbUdBVz
LTBQ+QMyyQfLzgyFABtpFAUxYVzxM5N4eN53W7WQBwcFsbIyXeFmhzJbHM6QTcgl
zYE09TnPMuEl0ylIpNzdZrdS7AlYatXmHIADuI2vUPq8CwyFxFI7McGb0UDvxGtx
l57OUzO7BjPL9U48ITJycz1+Yyn9wdrAfY1YBVdU+066eEYCEED7SjkBoeQShcB3
U5x3klGxtU9aMCJ/b00j0lYpTXcykt+zL53n5g/QzC/Eh5tVQO5Odtfuw0RaACcl
19lcKzZU2PYzTfx5DG1YJyfCaXNA55ODhNGb+4Pt7vUyTBSHBZCxjPre9td7AbS7
o3p14DKh5hTvdtQwOqdJcOI7XD+xH9EuZkdN+9gqcKieXWESLFcEXM/ZOejiMSR1
w8k+vjXa2XPzQmfp/yB1hemHxuwROELt6sg8zwQvD7jODyhH915pDNOIfVI6mX2k
eQKZuXfqMDnuDehafx1FbwhZrwVWtJoaDC3oIz7xKSQ+bR2pcNKgoZA++Uf0TZa5
s9NT2moKOGxNdTirx/WB/LWt+q2h3gJP5Lz6iCYt3nEDidO0hSA6j0pKg1uvBAiI
B9xVmqPScqjKODTTZOslyQaLL2ET0Sc+3KqLJHmQkTOd2HgUj9R8XAHMx992FGrB
FWt6UabObOIym1a483toSVAFPV0qjqONMN2TGESTLItN3tqaqJRgvyMdkGw/+HrS
0HtSa4lJtSnf4g8Mlnay6K4bJASCidhpqnaszg11pvCiY9YXIExZR1q7UGVWpIh4
aUfNR6fDhlMu6yJ8kU0f9c9dX6OZT5TdxLdYciIqiJl3BK4Ly1fhMzmZo/FLPiVJ
lfAqO6Tz3vGw647TCmTtSNwZxipk7ZhVbeF9LuRf5aBEhUTUb1fV29ip8dxiY0uR
CuYpCoCAEHo49HWF11f6TW2hexxHPX8nTvXhBv6DC0D1rxTBHWO6LgCb2FmntUJD
ta7ZdZYk0yq/N1pyNSR4jHCGFxsftuFJsu2pFBM0GtlTooRhPKD8g+j3ZvaWSsZR
KUb3I6vpZ4siV2tqkGZzRRU/vRaWZ4sIyUy/LRLCrwMxS4jPT//ZZcff44sjyOfs
YlAoz91eeES/NI0p+2ia/1wYMAeZ7KHiEZG3CEBmWyQBmJDttSvczK1ShP3t1QDI
6rnTBGVhUKLf8wDr4suHClTo6xJAvxPz+d6eu9W0R3VbUPXpzQH1f5i1/8eL/5BT
STkUe5gTfALj7HErPC4r9KwCFais0P0LlOQtWwlJcWePNR3hKox0Ic32YA/Gl2+H
uDBF4ISpYUCGFk3sINcAQWzFasmFx7mwf9v5x/4rKd2VD1bKzfJlQWBZZitLibd8
RKahtzIyz2xBZwGyS+omxU6f78cEqShIgkQezvWfxpXVr+g1RRjIUhlI2J5I7LC4
34qSCbvE3PTF+JZC3eR0wIAaphoHGDhEtdDc4pDRQhg7mOu8AKTT5/2a/vHRj1Wc
8oCyrbvrQD4rDnO28Did03RgI09iXX8gvI/GmgLfmXED/y4d6IMtKfittKlq5rms
3BA6Bq51VTc5IwhqJPb605JK5+JmdlSoTIJ24Pd13ked9x35R/jcoEDqpURuqxSE
j7psxipNyc3el5StBTjh2F8M0Xi6hMDqpsX0eNnHJX+JSeQNosnKK0Qh9fJdnZ7Q
9hYAREC4cy7N9xfDE3OY0TtKcTq3jOz+s8ezdWgmqWCxa6bWK9Bt/4arg9hmFmgN
/K4ww0SvrX1cWfZkAxxi+nowJXAf08y3+I8dvnpuKyhSJtl8LberAUAYc65rB1ZZ
EFNE3vobc3dDVAYbQMYorndFld1GTBS1zHHvcGo4lRSr0yo8gNhSc53OYgCHJJnQ
Ot9QKu1R7kL+pfIov6NokA/odiZPr/gWLOgxScaqbVd0GaTGDbQrf5AGPN8ZDtTm
PMZ0IDQcgUtinVlZ2GZcgUqKkV/UxLeF3E2bHT/U3vyjISOGyQSYcO+7mg+oOkGZ
+Lh6D8gfAfsHcTNS3MjwFpQoDa00WzI0N76pm78QIMCF39H+Xxmjux2DHe9E4uwS
BuIypDFyWCR8OyMmNW6IecFELPqzY9xWG2ApMcWToD0D48sDy5e8Xewep0SffhAy
7yvNQYz9/Kpucy/6da2kz1Hb1sy/p5GKYqUw965k3f2Asn55lEkZ6RVD8MZPsz1q
7+FaB1LXY5cZ9YZ8XIZzO8dh9T6+5yrtHCZ1no9wthWFjDPBVM5xQQdhlhzXBS85
wAoid+zsSx8WmloEuig3zfoWj8AaLJ4euBQq3cJtZbEmzUMS/BnZxmYYsiQ9/GNd
P+i8xvVOxqYplvrzJArz01jbyk8EwQ0EYeg9jbMVSKfTKKlpzUrU2P7ol8iJm20z
kH8xvjK6+hc50De7oYgMj3hAGCSV2HkGnFUmIFwvPLeUeJPDY3ctBNzxN6MbygRm
P1mD55qcvTza6xGpS2kFrbnGMpnGsTdneEU5CPDySS0041nMigUxo1J+wlExSL2K
0G0npU/La/X2DKHONzOZvApL171NdWKoZKgkVOVCPm2wgtC6sx+sg6dxEHMv5Nl2
LJlnvHOVe3OuOS7Chj8VAHmATbvzVWZXFNrWJaRrtDUyx+kuUFgHQktGYELwsgdA
XpoVbjvQixOrInxr5UzOW9DGoxY2VgrylyqzFnqniy+JvwbFD1LxR/d/P2uwk/Fe
1Nk+nzPCE3mkfuefwsS5Pn0hHhpz21bn8reuZ8uPSqy7Ba84Kz4pNtz0fdIGYxnN
rjMXKCvQD342NLseHHuSh0WflPKEAe2lt4s66Iamhtf/EFfaTC9uw/bOooheR3wt
pRclB9aFGuuaPrmdwVNTxBoxgifRNYKxJKH+dt91k1/Q1w7YF2mmWYueWUFahxDt
Nt+Ux/1Peab0H/zVR1FpA0+7us0FR+u0mPEk3EixBWmGUmGruZ2wm+GutW5SbfyN
Cqeiinfs/VF5VsUArXAnSqmEHGrl71STO87j6aM8jHIqJquGF6OSpsa9mhRWQlNt
uzqCFgwFWsysQw/D+AIEr3T1OWFA2OsDdpKpXlLKENaRzNl3VeN0SAUc8hhIWKYy
h+sLIJz+yikYsOHxHTPagY/IoVpbCmgiXW+QH7PQQ9IUhxcz4zagtiA6N9oRxqod
p9Bsg69UzV4c4XyXv+/d/h/oCdT1ot/gqVeEsPoyF3SD8/aW6wLOy2fypQsOsGXN
ITgVW7eScF9wirk4Tbz3qkumm/znYSRxqqEkslVY8LuY7dMog0MsUxeLqcVq2/N/
cs5qg7CWzkUl0p3eWRALfCbF2YZ45fgLxfiOzDGW8JqvvyoYXGhB9g6WZ5Ml1tFy
2P+3q/LWZmPUmhLCrQVLikkWzdep6tkmVDv0ej2fDhLU+YATCAlegO3slJUFh4OT
XPV6PoarAZYijj6u4tXuc0KQov5zrBktCIQ4hV/PK5iuPju617zYP8Z3p94KG+i2
kykLdrjo6iJl7s2n9bHbH0e6zcXriNIUAtalRB1EAz9WtR/Hy38L9CTklSBjpINR
PyRQexOrzFM+eKefyWMhOMoS90RK0RAGfMaOwxvclI4IcfZL2X3jdj47W/kVZOSx
ZkNnKAINoFLLZDCAPuQWh6Ltq6SfrS8VQ4DxpJ8p6jZGsq7PWKjRJcymU5NuDuwi
aKNQEAiTk0RjS/a1hbGP0ZL+0j7IoUpW/+TPwctvbn8hC2O6cLQF83npmZfBnetq
Nl4kpB9CbUXYcxCznQBN/uyAq14rZmHUqcuI59oSpaj1C7iHXMzXHiAoYu0FRLFi
YKhCU9FT4zXBwW5dzWUs15h9dBdRI2icETkA8uNL1cohoJk11lpSiEyvuWVLygRk
uRLTjMItuq/0KrPgrxH/Sd09LX1EDTqPfLAj7E64Fv4h43y8walKp4WDs7ibTFHd
G0t6lseOVRYQ8X17L5ua0M6PNeEydeADCjp5A2MVLcxMzvQhVzY+dpGyqyOAR0cB
hUtDiDAwlwbCHxFTpSaLgDgPkeCRkFoaI7hslT+TNXqM8wnScwNLYjLAdrrgiOo7
BbIkGtsHdHcJ1domjywVqRo3cJJXM+GgNhsKHXlhhfZ5coSwDggVqmKjnC/GZ+eA
OHpzDJAwkc/Py70GKByLkS1r6xgBICBP83Kaxmqr3/9suhNEqQUZL6UhRKk9u3pT
wwo21FN58pUGJ3EEIolAtoOJE8LfU5i1jba6u6T6OHob7kaEPUYlhAp4Lr6Q8Zot
eTz2Dv+SJQ7/zzLDtyX5gSnUHrQxM2UPj79nQfEYSOHtL7jVIN+qiJaPa+9LmVSh
3GTp91pFtXXZhk2mvlSF7mzdb2dO5yJ8Tjt0tL4TYzpHvLSFLUHeYyfeGeDvpxPc
wfcNQ1fpOAeiSKAMr5EfFGjh+rjm6TTtHGDUr8cOy75PMEU3AHdo7ibQeRbCf7kV
Ov02yOPzUgPuXCb9GP/RHV4kQaj4wXklyeBPozJLWZrs8vOJirQtYGuGc52UK9lm
hM4p/ojkaZ7tKDq6mhELJ1Avpm9K03JTqsfGv81lYh9iT9jz1s5jWBH3nMxapdpK
M/Gy0HKfSBBE1xEj/b8aUaFcvWQv5G8MOsa1CFKuZ+VjWDcgQqu8UWuPJsBzC8w+
FORecyiQ69HjhWOZtDmuhjBQsULlHwhe6mAYIouGc4VqOGHtfRlnmfy03uibhryD
rg9xTjPd6jkJAymNNIgUoFiIMYpxUuSioSCMQyDr7L7K1ybh2S1pDLfEf3xUhUGg
YsJ3Ry81AxwnrrjNdhTbp+ca2HVDfXHxnFWZ6OGPpPNcz+OlNokodT7oFr2lDCg+
OAlBYpvB4WyGT0pPXIgDF+c0QK7Yob1MpTtG0ZjcytvIe32u8rjBkx6H57HpxaQU
Ja1zanIKHAIQEmgvVOXKjuGRzoTxM05WiMhl6ECydWjPhkpD7gO+uz50A6+0Y6UL
MJMlWOqrkOGMKvp3WuETeqCkpUm/a20ymJMT4/GAUfZH2n5dOhhI2Zcb/xI3PcRE
0obSn+YeTzm9zUPXl0VQBNREm0QG1bn+kgIiOFQf1Me9wbpcbGdK7CLFpRhPwm+7
+iYRunRc5LkE35013PRPL5CwCmGc7wKrKKitJxFu1VJPcD0FvhsE+7GdItygS1nT
NuIk31fCeDZ17mL4IDXnxMGiIvWEDtH3YQy/uHDv6sbr+skwKOqi10thGDKfm5J1
WtERNa2owAFjK1bMoqQps1gcYJmQJYWXYQfiXszLcWixB2dEH3KYD+etcBwrLeiX
8BInf3XYyrqzDung6yv4woH8AJOCNPAUIgVY2Y0TDpQdX0bZIpNUXxchT3MTT/yL
IctIIJcTgK/AvdSRzp3Nrm0v6lInQAevtGnzqg7nU495+scgb/PQgdSN/5XqaOcj
SJDyZBykwdvRwgoN+VM1WundFKuUX5dFiWbLnj91C+iebuD6xe7JI0bsG5DYWvs1
7FttAOTpH6wbn28zuAKCAVDCO9CBnDtOzOTsMGoibkIasKohUwsTYI3ieueKSxJ6
1dD80VeY/vkDk+AGXtWty3oIPcDSfHktsjbnhegku2RJ4Wn5ybXW3K3WivAzuM2p
faBJm2P5JqW9tG2ZXEQDCkvZjV7j4qYrK+TwMn6EgdjXqUkZ7q9NdQ+AQP111jHU
/nfnDBsrVcqAhJvEXkTUvU9+9zn+vXwbg2koxsRy35TrLzPG2V4OtKOPj2gH1Vy/
uf5s8eJ6JD9aojcFp57+Kngmy1WCqoKjzQ9RexCUNby56m8RzWyaqyWYRJhY+/LS
ar/PtqWUmnhgKtHxa9iN4ehaLISOU6wvYuFhDx7VlgelS40uzxrW4DFqOuTIXRY8
Ur/clJiaZVVUQNQSlpz9DehvDMAuIRF3x4Cb9+FdjF1x9JAu9oalCpn442mrQ2az
qkArGiux39k+rk+6w1LpcrIDicHm46z7GbV1vnqkEpaA+RZ3RygrkIh6bSwyHXwe
n7O0RcbeG9uLWJbyVZnmmKCVYdcvCXtFi0WmKrT3IOeHCONKilqwqOoF5khekHFJ
pZnEKMzehC1OBJdQOplm+fmFR5Lj0awiG4Y7a9V3lpu6VFhpLB7X7evjKHP0OLBs
vAq6Onyjoz0snbzA6B4j7N+j+1b9gdlqZvZXnDqZhQ5M6fHmdHhuD1YKnF0lMgka
dXDQhf3/1nZJ5eKj/O0Fz9LR6UV0iaG4ki1nd60WYfPRAqABoMCa07O7IaTKM9t9
fhWHtNE4xp9mISKXn3ta3bk2eFwZeSVRBffqCEJ79/mwZ9Rye0UkTpcYe0IidtOy
+pHfuoM40KaYrdmngTaoUicMlj9N9b0ah4aeHmKaTCXnKdPwHh8vKQZ8gA50xTOP
zFw1LRfdOqQ6lutCilSbXZH5ioqFAcHo1BwdeMOh5AZDkbXzvpk1mq7eGSaSOEjZ
qyO386ZrDPGp1HENBV+9GlmbbDG0ltgi3Xy/zXgS2M8P0vOLB8qmQfBGkacoTbvO
pyet9rO0ofx1BSTg+Cd/vN+SO0HQNc5HM444aY75UT0Nl9eiFtYtmgrRwGWontoq
2FH+PNUaiery6Ue+x2rFOpH7IgsR/UX66fqrFjsXGovVUbLXcfAzCd4LG7A/DNzj
j2DjYC0VwHsk1RYD9YT7UfobQ8xkpbYQbft1t/P3QYtzQr6fWaXgsVdHXjSwJCME
l0J8Uf9AsGuIoiwRsokj80paa0D7Q2L+WThAPVmRtOHIc66jX/J94uOst50TO5yN
0bYFB4vsk4DXt02Y6VGURjHkQVTU9i/ym1fHEKZm1uN/Q7ywGTV14tT734Kvl1lN
YSZXOiu+qRqQz5bQwdkqxwHb9OMmNNpyZnsc+MPOoxo11egZQ1FkO48jUco1lucH
w25zMcroYTZ9DiDvBxpgBqD/2DuAZR3L0WCahvqe35g2H23KUj4UFWMhhF1m4LRH
fF8ce0vJRoT2ziorai23P1lxcD+G2hv8uBVadHKYTDjzak/dyqqbpwM+9x9X5ogX
m83MlKjECeKQP9ehU3IFn/CmWuDVQrp41i/TOm0dkahPt8v274Mi0mWrkGtaV5be
OT5qI1VWJ63gj07NVD+2a6wgd5OGinoL6mQnbz+Wq5L1HCqmIQwZkFy8tkuNSxMk
n3Bhigj0qT0dPvs4jmBLNcIF2i+pVs2z4j/EVUKZkYawjZ+1R6Y0uvtzTLMR33Hr
NUI1Pb+ClkXCgOQGOZdUCwZWFDrOC0rocImIDKYu9XqIYStcacyU2EVtdz7wV/tp
gednkuBK+EEijqYZnSUskYvn9IRtOR/FCoKtY0/HK9cBi/VihZ5i+8VbIAnEV4vn
mAO6IlwUoQq9i3uGQhpgmq8/i8TJNS8JyA1x0DiALFKwsTRWvkZPy72CE4zgbKXf
RoKo6jfAS1OG4Zikt7pGM/s6r6QaHV2nIsAn6RaOv8ykH/kimJDpyWGhomz1zD1O
1p/4Exho9r34vzFH+MW7Qwpg6YsiN1Q0VOuI9ZzdEfr1TpaK9BWBjbsQQWWNT8aM
sH14bRpf9LV253T4tG/hIRzCQXAEWtu+Sal3v90AoZMISYGf7+FS6xzzk1hSS5uz
DVfQ61vz+diPmMEh0p1VkaSIPIUqMmgTjb+xvHlefuJxoPdJRhJXxxXGcaGBz05j
ac/64iG/AHjqnAwOpNmYbUJ6hChNQvvw939/8nsILMnWbhaFMJEqmTBVyEX8K5Vr
+BIZFJB6hdzuVxvLmwug3KyoFxLfz6w9ViNPH5pn+7bj7jNDuoegVuccbCdeqCIH
uUENujX87gtIp36D/CmRhv4eZcfPmxD7bfrgFJaP+6WuqvesvHwxz5htuqUk89Yc
e1RjupcAG8dJltp+HtOYE2vjCzBUMej84is7EDzQ+gwaVM4t3eslqGLYb73AIcKo
J5lFF00gXdacHVkvW7pQNiOUQ2vY82vGCaXGkLtf2bstYDWlFsKw01tqwf4zlje/
U5hoPvMPrYbfXuwUT0wOb9QH6+MXCKotvohD/2Y2dl5ntVsofVIfWA/fuLDhyW3n
aJTVT2BjW0Wam3KEkcp2CHDj0+ECbqdG82QBAN4vGQrMN10ozA+Bqn1v8gFqtCFa
HozDoOnykkNaiUQtUkCuxTlvdi/m9iSksk2lRNRDxUMkQLZPAH14myv/4zslzKQy
a2RY99V5NQJi9bbW9A7JmL8+UNemu80hArzu4L647KXmsU51xtEmUPGoaly2Ss1a
apP3Pnld1JOiQuzyNvQD+Pqi6mpIn9R1akCOsWxALw70baq3EwLohPuQ27h8IgCC
C5pNb5SfUb61QHHxbW+VTjvt9smPCcOtP+NXFWB114x2cXLG14FYHEp6ojDk/l3c
hObRP/GmM1B2LMcCQMRzN972SHBtHENKUtWiwfs5JO9xc4rpYkev2Me4OG+V6K9N
ydj0MB51OZiAJJ7XSkVbSCtnNlNspg8EL0OHeLdDC2az4BvzusgOYWI9ktdVfxqb
ePTjy94Gad9SCM83/ndCmqC8voKQol6CIFSez3PJTyELCQEoVPqKNjB6kQDSa3+A
nxKoEkR+Uv49xAKv3misUhPeMkpHlTfkXFcaIxa6ac20bgus/BB9oTW5/0JLnnJq
CgoYGLSd76hXwK0kyJGomtgG8ludBwobVYaotIXkD/gdH38TYkd5Cj4PRQ6ZdatJ
QTcGhPSyOsmteMp2TZjiiXNeBpp94K03PaC/WGmLitv7zBnqUT6iWcejzy2MTn9m
CCGEumtEr5v0DZbbtIf7qfNwS8d2tLpp4BPScV/kJgWT3kIGy61SshkkzVFoNiAa
7cut6XC9+rDY4XpoABGOX6CgGXqHy1ETNBj3NTil6PyT/03WJUP9FRQZpS55pJxu
TCmOQPeLBIiKUxrBLl1zOkiiKjEBFfYiJamM7pd8No8VprmM9bMT8lMjzA2ztNFE
1bIrnP4MfhzlhgdmCKaZ2L+1yXvEPUie+mNoXdyFDAHlDOlF5r1VZOYkC8qfmiGi
d6FgzZ89LPASUvvr/b3lDNnQsA4zipSsz74zXqdt4SiT75qnKkNSHLOf9cSfMjdv
MxdQ82tO5krHFiwvFvIlDeVibJQHYjTJeZaTEW/M4ZSe7CAbjZKDKpEhgtp/v/ds
6tk2toGh880wT1r/61Pcz1dczOMYJbG82s6NFkBVxeEqQfvN+rH2LOp1v7OJWdCz
9UiO+g8Wpv61XR3WCyWz9xDpvI+u3GFGdbG50r9f5JRuqqDXMs9yO8ZkPDdx9uH1
xrObUEFZmuyGv4H0H5WkRNdtmw/j9WcsH2p5LdPXCRt0OQfOYG94mP85cUlk8i0y
br1rO2oK0FoqruqoRgW5v+DfA82u4/aQSKQmaUFg5E6Xot+fu0Vt/Ct/euTcERmn
zKfvUUZqT7Pbv0bEpEw3bjVaiCuNkbuUQh/6YSKfMziP1BcOoyDuGKJtmUVSAeoj
5m3VAGtHMgiVp1royJLTMQ6b1Lgq4DzVc7iuR4kenAyeioC9G160DQPg+SIEPcux
0McmpqfaJSRrQJ8CqqE5RShRMQw8st5e7Hr3huFquzkyecuwG9HgvJlyK/Q0XtdJ
zwFKcQKco3fa6UbR2ue96wQ7rlLhrcHJLTejPgg+OmI64/a7RZ2fsHiMF/JCTdqk
UKLDVVV0/B6CKbelh0KS7xNhy7+lhRgyoBApeh88kgQg9qw0RbRqp+sjYl8RtkCg
UtkL/A72TrLiJKza8HlPtiJ8AzaHTi83aVcwnqoddhha1Q7oYhPP37U/1Np5P2r/
b8RbjGYV0HYlue1LXvOIwxxeZ7HrTUlax5Vz76sMJXd2VQM5RnPDeRzrWQDG1Ux5
tpVOwjWzyi1uJLWowa5R9G+9uUUsa2BGs1X9VGiRDEuSgvy5Fg3Wd+W/nG/UWrJa
lQdxe1hxJca/U/fiU8W0ahuJ4n+B5KZFCHVHaDqaGHxk6rG0Hm2Ca0vmZlPvsmuk
83MPsZ5onY5HyFIgUyarGYBV5YPYOaPywbZ6VRHuPpjLtJSKrnTEXc/fVPP447N+
gO5Em4JsMaJh4diR05s+Lxvk8BdfboPZvm/oRAHdVj4EZO/wzqXbWzV40CweSExj
U5m62eljlJEc0WHGJYj5jTEsYW6GWSs/XhjZ2V/K+2AAgr26YBN2SALw9Z1zPD0p
1a/ruLIeZ635hLZLG892farsOn8/zESI1ltV9NBbXh1AC83VnuW0aMwcfx7m/fEi
NEoZLW7dsqKPdd6YbpulfNYtavYFeh1e8CaeO3diHAuKDG3AQCH7XsfyQUouKFd2
IkhPNkbsJC2beian+tmJd3+lbBX6Ef/t4ZSOoMRvtUqgMG+11vT9cj12zNkzyI9z
UyKkYiWgby+1Nc3xghPtmxVvb2/mWbLIFDAxO7liUXH0e/KyPFpkEBV9M6vTo4zY
JXj88kB0WiYcMx85Ce26g3BoDIIYNiYAbQ4dADFx3Pna0NeDmBBI6/Es9d4bW2f4
lDBYei5ZkWu4nV5S528dLSOycARaG0YMDsu4e9jnVr9zbxwpFxFejdUdBev/LFmk
Z1kxoZJql0EzSJCa3iartOYLzjbozkUcdDlgwqVxbcLUv6ES5l3fN/tOJZtWv5jB
SKCu77LyvvIZdVum8QrV2d/jUi8X9vwfx+BUnIq0G/jjPY/yNGtlsT9TWzBDsrWC
nU2f7Iij6XdkPIO5hUeaN/9X9NJrzw6lbfefevnYx62gc+uSZaEqv07ipsLyEDyN
/juKVWTRrlCzYxtM/bxp81i81C/o3dHzD9dIYXWg3r1AddCyQG4omzhtTnznB6dj
ZUPVt7T1ikaQALjaCEeox7I85mxkePb0f/r+h2BtgPTDGr3sdE8/RF6Z1xJdP/mY
7BNnJg2joAre3GB2ROI0mREm2s87tt8b6fQR8A8ljCqoiSYUBoaTFLSjF6nvw0Qz
cMAF0fT9qx2MxCXSMhh93M6pa8nJ1u1hqjwQtuEn/Q2mWT+gm6kwHM72rJ1dxMtt
rydrATuJfMEtfDGY70v/R0gPgGM2xLTnlgpfAdC1cC1P7oBm4AxS/z4ZNRE3/7Rs
whfXoM8t7zSN4YGydvBU7T8QiV9POs5DA7W3rs0vxYzG46cw1bwxdvSVq1MgYYs2
Tpup1U4QivZmKSwu3+bmYUap+osFqZzJXvOrULMcMOzVcUhplFSpbIdE+BokfElf
zn360qwwvgyf6QsQhnZfcyo4m14vAmtN8HMFdfk35P1JXQz4HAU1YFlT4hY/DNN5
OACvVS8ERDdQYueDqB503zxtj0OWikHon5JV8jSCFN/UKGz8dvTcAH6mP60eLITN
ZxFyuM/XiMQCarWszFDQWC4KPew5B1X5tOqcHWmubh6jZHKahrESRzCZ6zuw1Lsr
W1Ml9LgIuZXLswJpA2jYP8K4rwlIf72+PEWhSU1zRBZdpIk9uRoaikjiURBu+6tb
N7QS0PYAuFekItdFcwdDRlWkv5qAHbfw4CvlfJcltu2tm82O4FFLtkbWdpzrtiLh
iDoE9kf7CpM0+F3XohqPKRFTvuZRiVpyDptsVTIeW9GKA0sOJN0MVWuIqf9/v1fH
ND/n8/Mpo+2696KnGiuvwY/8x9E22WlAn2uEUk7jUmQV5u1BkwnyS9IBMgz5pN39
D4CEheqCJdfV5xKX12Z2OSgjXct+vgZY6KAgx5NQMAHOJYGQ8g+r9AWJ1Jxgnsi1
mnIwUZbRS61xuw0Qn3WAfG5oUUXEwQ5Ej3LgLLzhpDyaNw8BxvtxoLb7wHwCqNs5
rzqSIUZuX75rJq9TEohXfXlsCgPTixyWcUoSMeyDp+OyMHaVBubK1KV4lSHDUCgN
kgLs7OUGAyuVRCApefo3eRbOdKtLmPpZeSCQRLDA3oIJUho8OsEucCUpUxIMo/kM
xb7/8vX1qdEXPiOzVNoVY8uAztsLDCE1sNPf8RU0Is+hkNzEea4YeNVAI89EkOdv
6Dm5C/8Gm3o8O1U2LRBOcQTyzaJpC1D0YUyWKN5/kYpRdyLZy44KfHB8OfJdchDn
Mmz8WtLcTYPlVuyqh+6ON0wu84bB+PUkVVqgjWQa8aOIogTQ85R2nB+z/EZVt8L3
r1yjC37D37l2mjJxtA9oGjJ7t6v9N30TASw6Y+ZzaUM0LNg6DuNmPabqZXFTtgtg
ViqVrFyKp2LxsnMM+1+sHYQbqEz2aDUO3pQKDY/wdQ+YHD/gb+Y+cfNmvQOiGRkk
BfiYASBCSuP6gbtg70Eez43JmepIo34MisMv29jri6dBp5m+plhfTlsmur+aOAmz
SRXwQvcnMJd5JXXZT83kGHqwQRRZKh452Pept8sT6a3wyKfdaBYOrl/ERPpmOTYA
d9CH27o2NvSxtZ9rDmt9cVj2Fw4qdG/VKQH3vmEb60tLivGmxydUT1BonFWlHV6D
mu77U93ziem+eMbtOOaogS5TbghIJV7xqdj4+uR2fkOeZy4dgJ2yo7obHnU7c9W9
qGtSkNcuu/kNN8YCZZWCeO0sUn4kIGPb/vPAondmmRThbZGZGVxhoKbE9M/gQa9y
lRJH7BBbCbMWcIj/R20OqL3H+93w8dKP7IrHeizHJMFHDZrqHI5B/Iwrh7tS0mFL
uu6Uz+JMORMK9sm/obioQhgGRheHN19ScfjuuNXBNc1AEiqYvWUE0yNtQK81Kak1
HMmi5YDjzLk9o7AqzFAmlctJo4c9JumZnxZ1753OKcJwZsGR6jE+6hhsRsYPqBY+
kremVHQOCxtSivAtr1dhNJfy0rn5x6xnJfzh9upURX2v2Ju/Ah9B2XPFQ1tv4vJP
RCJW0eDIyUFir/c9aI28JdQpzc/LdnB1fgOzv4guRy5b4nPM+R0YK04zB/cW7y8s
dSTYXdgIQ9PMKthe7f5PcXmaQO8qI9VGpGxkP34lgbyriJqbc0ykqLqBT5hoCITb
Irj7MmELhN7h7lHyVHK0xz9A+fGycFnaR+lxMH1035XarQGWPTXEMvrPsLslfZX8
7D+VHeB4gGlu6eUIZ/TNsbtgjtE4YY8OnK3RNXBAayKfjHi81AJfqeM8Fp3UmenF
U6mlZ2kSL+D5lbqv5UNXxSkO+zVKxQEBZRUnoq8zwejrDofVZE+HjkHuxg09QwcE
wdjz9aTPAb0uxvfMXV4c20IGWshmV7rqhAIJonsAmbQVT40+yer6AAQaIZJQTawl
16mffV9sifOqOzW77JgW2H1/kBBC8CXi/mfQXcZqtHIy8/vlP9FzYHNXL4g5U/jG
q8bzeNrU4FkzJMOiUyxW9ax9VuzCfcrPzcfCp+BxddZa3bsg3m6uvuaZReGCIMyH
IdDh9WLzow7A7O1Ly977hWoaaG4jYmo+q6fbIEwV/mhdRK7xFJfIJWijrXdlUE5j
FBOO3q3Dh9BPabaCu65x8nSV20mYkYRIv/X3M+pHfym0acwLO5MLyqUJ580PysXx
l9X4b4lqi98ClxbNIuEERm59JwSOHXRN7TQ+26xNP8fRSX3fOB4LxdsV6lqXX5Y3
lEDroqPrzFHUmpruWfExWGu4dltDTwTzKb23mIFoxYCNBCM7+SB0LVDM3SqAS+Jr
fDyxgq0UUd/G5IFSG08zLWSDiR7YgjtJ19k71JA/eTwRPfxanFMo+bmKIHCx01+p
qoR7EzKZKRKxVDdAp2CPqQXzUydLgMxa3A3G9F9pxMUd4qV9IgksEuGggdeCGhjB
b1b8V9UV8m7Bid9n2X5v+lYJtomeA2mHBW6kOXuBw0XToe9TfQyTlIzZKcVNoaI1
jMlWv2m1Kba7f7HNxYDAinkevkNiVDjVYSFgzpijeEWLrq78+Ijrys4UiixrJ2XQ
KRpIV2f/EnmxqAzFW/WV/yz0dVCExxGLVb7dSWw2wgUM3BavwrmQdFB2KmEMLgUA
kvbjHX8RDMQM6ImmIfVeRw1Izn0fEjhHrb5esZ74EB39sgKhfpX/6dLzLizAPoYC
AMvhb8fWNbLt86JRBuidNsFlpUMOxqhguPcsRNaOwxZ6hPxxehBmq8YmPTikKoiU
MMJVsfhpGAxT4WkVTe0fObyfqAHmKBmMDACk53cQhWMH2Ai4qAcf7MZuo/RuEx3u
3FFAJjxX5SdHqPv1lDPuLTjqDxujzkDcfeiiJjZxlj4dllAX+LU3rTqQhFOxUnC/
LWlRfnLcBPLvRhku1Pk6wK06qy2+XO6S9L3L2h3+xdbup9g5wAO+C7Go/Pt1gEhl
Gk/xHREqjW9lOrUQxmIKTRtXSSp81zdcowlMWIOIlTx8jt+xkF5QOAp7GkomaURV
bBxOpdtJChVDphzAMIaJMe6EpHWNwygpkFTSVAfyjG3bouOaqI+P2tnaD5HvzPy2
jph/K5XeEPqexvLaDVASio9LG6U4Blj6ClHHrlH5MuxSPxgorfGGGvSgCgGOmnhS
PyZGeyW4OyLk4rLtMyxsCHYPhqHgSGS/CioN8q1P6+QwEstirnvN0gJqaQXx3zf9
MksbFdSCNRW56LcczIdJttXmD5dz+1x77qby6A20ZoQcSWbNrxzPSEp8orRPG3tm
PLQZ+YEfeoqTmwC9KszJMASogedc7XZ7a0jv8Wc8xNvS3NsTWuFyfWltfiwsuokX
R9P6IiJHiWPqfTu6iPThHhDZCgCG6rGtSj2t2ePNm1cNFlZo6Gh94y3XiUSmQ6ne
nW57EuH6uZKsGmjnf+dpSRSLd4EQPLoTJ51Y5eycj7/Jg7a5ZdcvaIGrbmgDfqOj
PskjobFlJpuMCSGdnu70wrlpmi6MypyBqV8g7rAdc8DjZWZJUxh/IU5/oQV7JB4t
UDB2iQeEkmE4KwhvbNF/sp0XB+nHEbr8FlUZzBvOSJoSqn6dKEhgV41xKzIEvnbO
hhJAVkBJCT7LEq0h4Vi6ce7q5vfJNvZGGvu4ZPXh3SwX2zhprovCOwN53guIms09
8Dz6abCdy+brOPVYIaP2RkZ7Rrm8erXiQYJFGFkrp/uv49mWAx2ZCu/s1Kuata7D
Lrro4hJ+E/+ZPFiQaTQKSrggjd91EpRpUvYY6mEeUXwuJHMTx3syJQU3TXO+YBlJ
nj8cvPrpzzoRQUdrbR3a2Xjgsxb/UFwWmolYxKNo6PiLU2lSvMj+8f2TF0T7V6YJ
2sk3VIqrY9kHnj8Kc9NSyynNQzc37r0esGs+2beQoHKS3b1//99qXdKBBxkK1+7N
aZwllZBAjN5E0d8zoSL4K0djIn2VGH89kuCIRnpbdT9GsN2BHiG2iTjJf7VKu5me
tznmZ9MXidA9vmrIvik7yvgvmfpwqe5jERzKsP/jfc4Hm8RBlm6OTzbLEdmAbTwQ
XcnNZFgUMssry0vZwaFM9dihb3mEe8tmu4rd/+WwB2bkp4hhJMEg65EQlMh9FZd6
OHLP/Rah8zsEyXYlHY957PR8yjIgEnjmbZVaonhKZ/kKJwIhlhHgYTi38ztD67Aj
f56mUc5yl26E+6Yaml7nPFC/ml9xXEWIm72HHG7RbHor0rsTptff8JEyavUyw2Ua
b43meKLJBQogoU30QTabHl9Xj0PwfLVG2sZ7r8yWsvzgWNoA4XArjFUyvfqbvWSR
cFCciJjp/RAM1Gr9JODJk3q3fDlf7u0inLDxbVc0rKiTGaTfHw0X6ENF+pOeP7Xv
KaBN16WNzdaDfNI8x5YqHtDlyec6drL7pWSj9U6OXdO5kPPEhE/DT/1ddH1w2zjo
TzIadOyb1fXqQKgzG0zhG9hP5HclMUdOdrFOIpTyNtVKbn+91+zEuOdRt8bcooPR
cAph+eXhUQA9LpJa3wVPSDbqpZ+rj/ZtYcNsL/kg4oU0oYk2nA720a6tXO4qB6v6
/b85cJOxl9hGQMTlOGvCqN5GXtk4xoYqscjqcSXNE+4ZMhPQIh6H0o4KqwgPDxjR
9faKHCi5UD1XN3+QNp1f1Ki7DPqpXuvVokUCIoPkPgAj1SWj6orHJQRvh0IREJOV
73wvAms4VMaxTJoZNttt7PvAof+kzT4nUGZkq5zZk2CWrmpHuojmogK21TYTedml
y9wISW9RorS532DObHVZ1JAcTjRxlZzOuN8shsUezObNtPCJzs1Fpu8BVsTEK+qW
MLW4kbIhbhfd5eiKeEr763gs+2z4Ey+1bPG6Ru6vkBsWSdmGqg6llpi9YmmZlxWf
FUuH6H0P2cU9s3SrOY/qGwhoOmDDkXyUixLoAU08Y+JR+syr6klhHLRRn+VkCHiN
c9tJZ5IbNm/VDys5lqMlufha7+F2t5Le2j9ZZCBB0hk5ybZDUXuvhhS2cUMDQCYT
SaF2YS8geh677ycpvKz3sEhiA6Cf8dHym0893XrVc5FQkYjCyuevXkqUv90HE3oq
0GtYXCIMh5Igp38wPURzzBhy9jTdTu4KnTEYfwRyRv8SIVwZ0IIcT6T8uvKPNzZC
GufF7YGNlmHM0Z/ItqZCDNDBuGj7nH02As0BUpobgEPp011+THroRpVaonRTIGf7
RNMX78Hu7yXSfQE6fp82E2qp5pKij0rVwkqKYMGmZTSyLR2ZDVMniCHPFQyOxIYW
S3x7oexDvgJxJu1RNOujPVxeKA+Kjx31NftMuFSHsFaMwBh8firw/buyxeWpP+2o
9yvxfIzuTJUhh2te4toqjpK8MeWsYWDywTxtAjy2FMjp8ODsMteb5gMOf5yoCri7
zIiWdIG7DpfYV0zbOT/F1mMLR9If4WTYUyHLQ/hjWJDcE0s9BANM3ORgVXWLP5TS
7fSty6bSs5rUEXuewZLqINemOWHLbWAHks8DbZy7AKpfl4IwUC8Vat3eO2B7bXsu
Wvrza8fdO+wgkng4hhRf8HxNrUnxSEKIQ01jp4yu2+XzwAOrYq+vvEp5q4dRoBla
zGclV1AwlcW4IumHI5BqoQWMlEHQqnAg+REAo9eIdqsXoHtxb/VmfD1P2SjIfgz7
TraTDzRcfS8gQZqWWlPp8AT/gWZYAX/lGWj7U7ExAZPGSnvUUXiI13XyoEvr8pRS
zUux1QMBLXh7jSxIK20iTsReP6X3dTDxTsPByRPlh/LhUYHK8Sbe90PAacckGFiv
nFIJ6+dVWqT+EQ9u7z3yAbUV7PbmAOIH79ZjonmODsGgUX+wpPkGePm7tZs4h8oq
H/PPDfKpOF0yBg5KJq6qk2ggnPOMmHweX10HhZbTvg7MyxD9nUjUnylsaeP+fBQv
k9WD7zg56bSRqco2cr4eMzYulfaeQ+OhA6NiO0UqLYvrAgTpmfDi7doCN25BmLbE
nxk5UZRce5unkGwnvrK+9SliO+DfsAyICWQXIdpYkUtl8zL5ixfUWqTWomfyxyoF
BGVSE6mwX5tODGnmaS4irCpgwdu0Srr7uMjOjA108x6yJGqZQFHgJggCtziL9IkZ
DnuaMHKxexKXzFPi8EVn5NLqPyOQzXc+lHL34QbtJQuvNyA0sFRU/gBTH0dy8E4l
LX44/k1aP8g7snn+XRS34HVRwrS2Pr5Rj9ni9gdBsVStWwslWLGhod2+lQfjg4rw
kDHUJnmMrCkFKGUPMtGJnmxJctOPLo0/rjQcWit+JGd7Pe965UUm9oZb0xyQE6jP
vjBwefmzMOgJP6zDemAXzWOAa+8om/pxa4fNqoo+Apmy9rEt4gy+tI6tnI6PpSqO
M1YpXTr+RzSVCGCBvXbv0piXp9mGZFTMOkoknHGtsnMULAyJikBQ8p4v5tVrbpum
GOk8W6iIrAKiF+jm6gzNkWaTiAhN+KtHLMwgY71tczfBJz8XjcEi+ErONHhyz9B5
By9m8dJSMiwVQRlLRwkeDOnDUh66hTdvQi5aduFLJSKaPE++V1luB4dAYiNwsekm
CMYW8DTD7FWK79g+pGt8scNODD3OvRoLB05utPlXGm3RIdFnXVp/Fbhjj3rPjCes
pMSWMnm8WBi2MAB6jyzuqUsMJMdDF6U5CMP28Q9hfopVGf7lGjv7QAwLGWc1Uwsc
MYxUupK8xJUbLX397KQ1cAALnSh0DN9irpxNPs/qU+StD5Hmz+Xs7+/DYdfNh0nZ
pIZa24MYJatY9w5mYAi2TsX7iJ8RucbXmm9V+lrlwH8KcNXHAIPEZi1RgZXTHCvH
7v+mVmAOlz7jQgh3EqbHMtEYL70j7XmRrOvEjJfVyq5rRJAxIeyPUbk/i5/iucp7
nZY181pYpON0kgpgnrCg8dOtp53Nq3zbmbQqDMJRpcZ5p0r/8b/ugiYSQmRg//4j
VHB6rwFhs8qUL3PwqPDDkSa5ntRMs8ADfXLSdUZa2tyuwR69SnCPjhyI65qw3ihS
ZpC0ryu5VEw/ecM9XC8O2s+ozUWriXDCyOdt1R8DQQvtV6XxldbtfM1DCTDnzdMO
rD7o6p96LG8B+MKZS1LZPxBki895h6k8DCnW4zUrJ6EyXOgb8Jr433qeAsoNYHok
6xaZb9veU9iPhtCdmc+PPEoHYMDr3tvBYa1f5K7YXzo6gItgsyW9ivy7v3h43SYl
CUK65OfNA4VUCWEQgVjXdDhykdQqe//PAC76tCyVeU4ZAqVSv/D7weAOwKWljQSl
Mh7W21mYhChZC0b5bKV9QzaxuxlIhxOI1AFme9XhEz5VZIfSugFTo3fGYkMU/i7k
U+z75fLkMKqRhxfejk5m9Qd/wusTt9FQBT7SvSmioQf8N5wS6tGX4SeFqgiRuUAX
6KKvEabF9EfC0YAJQULzf2/0LAH9gFmPCZ754J0SbHzz4aWvGPEV3+0rgB8+tmkp
SYn3v/zXgK/KIV7tc0K57o/eLuu2ku18f63skJb846VZKbTNF9bpJS5X/0AofCW4
FZGrp0aet3u7PmYCHrDLFsK5AlzNBNgHLwC8htBKWHeVSHZ+TBhYRhkD2YIkcwaP
ESmnz6N8Drm4ytBSXT9aZBoqUii7Xcpdaa8epeR6V0NDDTvSzlPKvPeDdokQeZQm
+eGBVpYy7CPePxd7PCq25XmigczYwXMNvt189H1w1a3gH27x5rVcShYktydvp0kE
omne6jSbQmzEW5v8tvlokVVxvPVji1jweE77DOExL8VS5qo+pPqcF5IS3XCMNoTA
A7hacO1X/pUif+hi4TTWirB72sG2LjbGi+sttRz27Yrm/l4PFv4bvy1wtXhGzBOL
8RADrA5HP+IZ2vXbJMVMz2wl2eEzRUv8E+iZ70dSwPvQR7FVN46BLvcRrgP5XYLV
4Zct2Luq8F/Ib8a3auub6Skt6+ZWmOX9eKj7mLZoYdTTQs7SsQbjDO/DmS731+gr
oHMxnqZCaZGdD85fFJh95zXDg0SWzcqTyJXCRwmHKSOZsVUKpxNhyRr37apcOXa7
BS61S7HPuUsNV4wvg9OR0USojThhG+hifPm9RB3RwS8YtRBwlqJFpmmlo5oZKYJF
L9383nsrSZ3c/5ls2B3glo7LKkRhpHe7SHIJFoqPrLDeNr1b/pPHA6jUvlGceI37
vC+N3ZWiCFX9Ip8Pa7GMGnEGCugdEJDMxU7heVlC+Zb40DWuMTeDi/Yaha3XewYK
Q8aSyrDaXNv2rjSxfJXEF9MAAvTTPLZ366duYeXltcFyDQP8ZGf5BYXxlIkolAEA
NBAT97C0GMHeV5s4BY9AMYUB5RiTvsYHwMO1kIC1dIk54QkC7DRnWQ0zaTQz4uo8
PVwZ+AGpPLnxpgOFyiALvCTE+HcdQCOPYNBLlAJqr+BQ+3kxfndqN3oIeMoAkIAa
BPtug7lsxwFfiUEnmzQZ6SJturGcX9tDOSr58zVSZ/+GSC9vJyirWRkCiNw7Napo
7O7vo23gEwjiU1XhX5/WW4HbYxvyFD8Qe6BTlezWxOZF4FH8onnXgysPXiSK3tNM
2JPN+c8gWZaZ5loNllxK1BxBJ41yDV58pBnQYjsYLuWp0B+57rCUpPqVT32hJ2aN
dsdTQSo/hWfpa6E4gWqKRG6UDo8FC6H8NIJDZPbiz2fgeRPySZVGGp06mTmaF6g3
LI/0JYu8PuPpjEG3lq8bKxjqgSK1TbOSNd36VobEovMu8IBbUEtX5FNyToq1gIuD
v/jOkpqtoYwpAsGX5019iPpOv/usUFhDGHwgxzQbiX7GttDJREeOX+hNmAhYhN6Z
Si79A+VLy/Nu3MBvjnl/j+5c4dbCVSYHTEYWit2f8T0zpC1IkeejJk5hNSoUBy80
OTjStf8YucnNoMAdU0fH1sKLq9qIzen1OLSgM+6M+OX7G7puj2Y65YK3oZXxWoky
hQ6mzzOi5AdBhP3sm1jR0XiNh2kJF50xXq5o5+W0EEk6R38CuZvs8wdku9+mV1NJ
BsxWzJ55Ae0Mv0wnn73d3ipDg+5GbAfbc3CSTnxV++0Gx+d0ODudYBnfgPOOGjvT
XOeSbhItEiOx3C0zyW1okfpPWqKAUEpafPeM73lHhTMCWycdg+KGP9QtqmqyTGkr
h4DdUXVWKSBeRb8Ba1QU3YZTIxT9YttenZCrcfLVg3OQgAew5ZdxyzekaQCq/hb1
loq/iBNQD/bMw6aJHl3dc0wH8T4aD6xPf/jnqBvbFitDHuU2ch7VACVYtNCDCa1j
5cXfGhoVyOrlm3HIHJPmQfPXjbXbl4IYQswOShWK/t46k5VRoNzRqGCNazgEfgwK
tAy6K8im+47s4g45Ntis6BdgHWlcvx6wcqfxwLwVi+ttItxLxRJ3hOFxa/T6beKT
Tx5jusizxZ21uGPUMwS/688gNqhIAMwLHvIvsE9hrUhpqfcvzztCWbPnq0GXdbQi
TTIHWcwiaklTAobxHv+306TMdncBpo0uE/0/2EOQ/48hRtZbEqBctL+aMZxIIYVv
L0mq03L0sWdzxQOsxYICOhVmheCSdp1ERfmwzEEGATElb1L1a05k/0xr36ZS7lBg
D1hnmAtHcYWacIfSQu+qM2bClif0gClAxTOWKowrQTXLy0F18vEQa6csqAYUCzPr
uy3qabiA+7DaqV8aIVWGmrY50m1tFrsZaUIoWFVEbu4TvdhWE/avVAi159zDeCUu
qgxpM84B8ZfntMC6mTCY3knHtOoHYk730RQQfzqOrgMWsP5ZGjMTUKLDk/VjrG1M
J/CPWMXc8w7eC8OAe1OhXvejG3FALJyvFOCgCLk96tIFUrVw8gSUCeSjMjXgiAFB
sOSNIpA4O6yL3PBVG0Xh3xgp0Uv8QCA9ydesXtiEKmkpwWZo5KujMXfahvpcew81
cvGXXbxO6edM9t9eV+aVsddibtszqL3PQtUo85Xwk/xXcTLzHr8dJorzvZwQD/A6
dPchizXyUIRcwTROoyDD92jabx0+EwRDc5tRVoOw8sqeqDRX+1OSj36xuTGOsz/M
tLspJdB/mS9ngegv6q2yDLEas+2yB6gcIN5pxM++8AvBB1L0FVj/ZlYsDZ1daXTC
q91dcqzf/qoNbI4GiVZkgVcfGLFg80FReRBMM3T4VtrLYcZ8vIwAWeZOJFsd+tRL
OVNXrP9kNBGcBsJM+QgUJkcczgalVVsBYCEo2WhPRJ7+kMa1gLyg1+mCCz9gQ9SZ
ZfhshL6di4VIjKUnm7SPWe8ihvWTvdFzyMaq81JbAZF0UuNriHz08M23CvWsmyh3
1hcHOTrII0J5EFVH5P0W1JUWdx5tf15pJqMX3dHgPnSZWDfAJutvi14D3CkdF7pg
RRUmjd0T8kztiF0u5ZoQAhbyhNBOTWlQ7MYZ4HyJFUCfP36HEWNaBh+KPmxEHLMi
IPL7eZRWPuEbukrtWmBdkkDa8Rn/cJu8dKbp+QIOIAYdXOWQemAMMWiBSyoaH/qQ
/cLWDc7mSoJiDzlqBh3mMjVUJZq5m8YyqO8gFkQNBU0knsKe9w/rl9aUEXnwCCbx
7uJj0msHFrzjFjiHjwFwzFsj5/pc3zg9HbdKpSF7CAxwGy782lE92s/WcxZn5l/6
eqSFcHaGxBxbvO5LfOgdGFTIYy5xbwFT9Pva5MAlQf8h+2Up140D9/lJTPEvWVca
z9x/13FG5DkFAcuc55gzchJlLfsHVj/RekPCeOdgv55xZQV+bj0eomkuUNNclEng
LGxEGEbt8thL9+86EvkYfOsDt+6KsYLz7KBIsfARfqz5m4VIOG+qmC1lcUUjGw/9
aNR1Ln2aqBHO5gIyCS7FIUNbOQjFglqqmXiB9Pz7CPJIpq2+JosNKnhBxvYhDsBj
cGj+5t5X/yZx7KXkhvyZT3yelPUej2MilPlLNXkx0q2zbWKbOlKkZYORCNKShXh3
ClLX+T2XYFMcApMWoVjKyYFd9/xQ52KVycC65RRKHzXc+7EdQdY5KW7Thkcq9FoN
LLizgSIJWzMyFcSEvezDO0vbIXeMCg2xnCmDdROahKwINZuscJz0qdWyWwG4ftrh
RNO7MlsTUmN57Q0F354X4S/Johb3iLnj9ArDNDtdaB0ryl2mflmE7QTnXj5eu/2z
IiNBmY1ZKwvmAocoqggndv3RVsSovC4xCmujqlxnT9jYIg7whgw52wJWUPlsA86b
6HY0qTCqSnEqiI9M+Sb4ZezACxY1f5vXWDBjFBUmF8V5SMZ6F6XAb3Z6wc5uzXgl
cNi6jCqVtsujRWht0p00NKAKBFfWncs/3ECuCviTJ9mMcGP4mFeZlYPWL66Mr/ZJ
o5Zh7qXzz9zyWc6yTOfiXy7yue4hYxFPhsQ9ZKyfhhuGbHJw8Inl7ZK8OKbEW6cs
xmyPnzmPsiYtGDLCtC1tZFms8HvjJk6LOCgepRFUKrnTmgdXMvGlXtpePA3D/arM
ph2jMWQCphOBcIQCBu23BQh3OUdvCmGL94BxX+MSh7Iycs+TnaqbH766NE2JaafB
4wCFnz1est0WyqxWqG7lY6dhBA/1GxfuAYJ0F1kdTlzk3rN65llAB5CiqfoHbgaE
pINr12PJLG6DgRRax6SNlEUi/9DpGYacJ1Arqz3LbhFeTBrysvjVgq0E+5Zdzv+J
FB3fFjA1aEMbE/1GFKrIqBuV53AZJtSJtmczGcORd0V1n15NhzYo9vcZvvs/YXfk
CG6xecNwk5xXpJn/DtM/7y1n19/uWC58UQwWa8xQ/SLciD419RSiY1yLo0K/H7bA
ziGul5g0EjK2Al53rw5GJ+oTOvS9ISt/4CEJ1wGuHokGKkUPrZgtgZPvmz2T8diM
qzoErPk6Wk8fYRI62reEtx+JhDPJsdDead7OoJzBrubuss/ZSNPFfab0YyVOevOh
iUXLQPudfcnWT88q8s0IDxgs0/QZYueJD7Ddnr+gewBLa+54yQL+2fAga+RsViBX
4yQ56g/7u1rXlAQLqlE/0RKVKWp5W+3AT7GTMqSqi7GExq5/RsEwg2+eKmhVd7S3
MEqK2KWqzoUAPLdTThNKVnJD5Uz6evADROirI1b47pbwyGM0Fwi6QH5oVH/uQntC
kszMcCNqePFQ2T4kGTgsVm/dWZGt+6pWoEUEylVAhig4VCvC/qRwj95FI5y/Z5t8
8L+NOD5ahKOxYmOCSbdiG2/DMliJHPDYD5OEvjEzYB9j1D2+xW6sqJ6K0v8wpZ5w
sC1ZJ+a8axOlZKUSJlXcaY2NZuWES4hBXrF4BO5uD9RMuPJnm4gjrBkewx2sIOJJ
im8nBujb6/C9YLfexzOx//qEwtDzK4B14gKBTB06kz3YFix0S2g1y9JasU3WrwEP
0q4fuZoGjWDNZFxFcQq9k+cRNPbqw7DmRp4DwZF7J6xqBLBf8JgZgbJrFjcmYKI5
Zm1QYASAXvd0aaSK6XFn7gj9RDhAhQvx3L/ARkuCDM8mq++QrNmkoxJCS89Dtw9n
cg/aNmW4IdEysHFhD+6Vu6vMZJbOdySLLbdl6pYhJ0CO7oGEXvUC4KN8RRF3GXwN
rnPWWFZqmZu9ATboNcZFs/qIDN/mvMW4cieftFP9mLXARUbNsRTBAb7zf8FOfpEo
B+FoNUiksV6hpvB3opNZp4ovsYZpWHdi4BHPXX49M2VIVDAkfL1ig2tZMGXYAWUH
rjjQfRQCv6iv/zbpHU21w6FVsK01qRFu47nw/hPxvt0vWv8WAMsWGU5wwOINUxK/
WAeM+E/Xsi4z2nHMKEVOhu6P64g1Ati8IxWZf6xvOB7HnNv5iFbpvIxFl9CDZ3Ic
9m8XKCiGmsD04bV0IBfvr7b8CohWUo5CCk6j7hnM/LHKwq1D1Vap0KkhxVo7e79/
h4J88MPlZB3OjgAiWFmRYJSB+o8zfFkDsb2dbEze+6Y1Eoc4TNSIdQ11CTHDyZHG
Re+uwQxctW60o/+t2YpupqJ/KeLLkgbKusCXyNfYYxydbcLtmSjop42J3d2OjW6I
ajjISqbwrHGh3wSg9rgcKIyLslOejNe/gSep2+3ppwFjJ7QfnYRodBaCsl7orDjl
yhZYLPB2BqV7C6OmbhiP7AFOGYQaVid3Ax4MYzyzzngZU/wtasAPPwrpazZkkaOL
HXiMewoxBOjADFdj0+pIGEiLQIMVhlPTgK6LRyqbTlaXz3p3klUD/gyzMJFD6Hrd
OMQ8dDsk9hrnFVQRHpu7wtKcATMCnGWqYX4on3/82FZF8rZft3vfSrnCA114ApLo
n+ghHQ9WV9/NMg5By04HFil+ly1Aba1t7fimb2GCAudFamkQZ0fxJzwifckhO5ep
j25aNmAOECGCG/6nmVIDuZDNcmDMa5WLzMYgBGCNWqSwoTcUCJrkI1v5fU1zO6Dc
rWk40DVRHeGRpNX28XhCwFx/hH+Ah8Em34Itmi3HcHtoWrUFGooudc1DDOxZKVYe
5S/J0GhN65nyzHjNsoWL+oem9gIA5jf0L+x6oFhMxtMY7vZGlTd4DXv5ET3IniAr
fWM0ntiLOJkcIIbNqQtroh5mTTkUi4M2+2Zfczzk1KPsKaqAM3T1qDmNirMmxJwL
R4ugmS9svTvnmhC+uttFpjVopECe5YPDh2Qy/e1yLFnAmIvseqf8i9ETbcS+NOLE
lu2+BYlgEdtmBp6OdNMgMpZLwQtwBYrRt9YqZQFGKPWJDm5B9c5Tcx102lLNsxzb
MnQvMmYNgM8618QxiUGNaTEj5TZnErIz/g5kphp/RAdvWWcNXYUMR4k8peDmCn48
Mv9QWiA4Jqe4cRrofTkCzyjTJDPOWJpP7oHZ6EPhaax8q3hKPr9y57maN5IMv+Bv
HQWzrdTo9ItaZTaGD6iYwM9Caz6Wd84YYi6jGyOXIQn1VGCLFSX2v2tsE0jpq9+b
kahlFwvNfHK7LJwasLSLVf8PJvdRGUywWiMlMxj0/gpnLHRlqC5Hjedh3FY0TNYB
E3QlOne7Q344wmXarDEaOQe87Pbie1SD7xxs/GeOF5JhMCL1B6mJsYntD6mLaoU0
sJcPhRatYVnmvdtGBWrQKNKqORSKyoU8aSRFUcZB28G2BDRSLfseHJiFP5/EAg9N
jf8iFgMD0eG/NpPJvmtpswS4OF0GvlectV9RhnZmm5gp/2TYKbuzLWNA3Lw2VGVG
L6sjIc3P0SsyKh65FW06JIs5hbT9EdA9K3lp2rhB67mFFU1Q2Nn28rw4BXbQlxjo
5fBcBQlh/3K4rMzxihqU/feDCxD+7fcFIH7kaevvP1PGx99eL5bQI0/UTaO5H4gu
GLqO2SOCs//NIz8AV/pxlaoDjAgUhcsV+hFauXm4uYac8+D2TpDU+puQwYMKe8KK
P9bR1r0VFLqhGDXsudvEX7NbPOynM3AKwICf0mHEQN6R1mB6Wogi2uWCNDphlHSW
B7g4pieNMqtY1/6uwjezpDT9+/+FsGRpI0nH6bk734wvOeg/S+x09OKiqMU/llzT
F1y4K5izv2UDid+zByUnujVxthNofyfoTs4gMCzkBDALUdUjENIJtRxo2krlp3N7
A72J398qxzSWVKCs0xheXUnwic0dx64XyWNkKLnSEP3LSMyDvgTum/q3UQyfPpH1
B6H9aKQUQTROcRGpuFhSOL5wK+M3kH2XrS4PhHGEUyhSdpvWCPjlLXOFkQ8QYQRL
Foac1sZNQW177dNkacMJZNA8PgITClX+qQ4mputF6ZvKmPPmxMKzI+WY+AXy/7iN
M2MkgIpQ+QYtpxPRPv5A0ZvXhXo76E+G/mD+/C5dtFRRoCpoYpS6N1Dd3tO/Ws/5
bQ5cpZj/Dz5XknODLUJb2VwNwdFxWrBWDGkY0jZV6O5PGEImr+RWedQJZo1IYrE+
mTE731dvLFKT50YxN+U39ieFXZJZbO0D3IMA+Gnq1Kh24tCjiy7W6IT9EL5KOec9
zjZUf/kgPXMTJMIYDfAw1pRi+e6m1MZsRAAeDAzvteYAwPer2VaNQVuKTjS248P9
3i96WGnAJ1L7qNgrMqPB5rEv37KD6FmnmdwEbHCZWVha6G77JA2BzgOO30/m6B42
lZ50rLRQ5OQPZx92E52SiSzPl/Dpbc3xQ4LF4Hb8a+4Fq9eLVUTZsuhGzMXD2m4Y
Sgjyzd7F7NzpwcS/n3+ej1Q1zGD7rxHFDSUnYvbwedJCLsZF/FxJ0/jW87pfX5rq
yF3svA3U5Iq/7QBIgkeNvpMqfMqu3TsLCUtEKUVs+AgQFPVWFUi2/A8/sJIYNsr8
/wvLliOh2QbblT5yDzjqNRmdYPkinzS5uv6Bp0CFh7t2Lr+v7s1eBijz4YymYLRj
Twemu/FXTF0xq0ppKfrEGPfeY/y6kglaFMGXI9JF5gewaDfc1tCDU8JZ9tnL+f/9
jGYQhs7DAZmHbTyqTDyDYxhZp9RYsjirFotaQf5jip1CJTlO1scfqb+dv8eKq8dG
Pjyvtve+0caKavVwlkpPLOVWOrzsjQKgp7G6y9qJP6Kj1mKdli41Ga39eyBdEtnz
zBBFOvPl8XiXX3Y3D5lAWlFkIvhhpH4LKefXuv8LmskxqUkxnnF9lTr5ynk823FP
pwkhOqG22s/9Bk5C3SG7CsSoPrV0Pp34paM22VeNG2i4q031B8mAjMRQcY6GzVx3
MBi39YUJl7MfmnLF2jSQiWaz9ruqc4yKI9ODriLI8nKyE8RAo9FXrMQXHByCkcpb
Qkx5R4Omh4AKS7lswO0bZo3Wjq55qMu0lJFm9CFq4Jhhwyp6QhWu722TOsBeGgFI
vAV8SiVGfbGATayY0ufiwjs31gK8DoFDAnAUf+HilQAnLEhaye4TtNZpZshMSyvz
4EJ5goU+m96RETRDbILDIekW/7zeKdb/XLAcXM0KbnnH59VYovM42RMS/NiMg43c
gTRyh29s7d4B8eA8+tEnsPzHK3u/HJTsrumcSWzcxV3E6Cz7Bmc4wrRyLZnPUJEC
fSWu2B3u6KuSITrm1V4W+w927Oa3cZbhiBwDfF/9xoaWX4tSuE68gP566bXGtRpu
LGtFTySXCDyk92xCoRMMj36jEFlfhnkiJPdsaVrTXekEkmWED0Wa71i3ytBIAmXu
BFa3ydC8OPjdbGZrrKCAP5pyq5q31RXS/Joe2EglqQE6dhMWUPSSlFAriOmjuFdk
721ubPXOxOBzYOu22RV0ze0Ej3tZ671S4jWm5+b6ARa1ugxPLx0fjk58Qh9PhAra
vQwJQ4TeJSxeizsvjwG2KFIbxrm248U/fk6hcksY52s/6ts0HEaxfT6c0oAU/+hO
g0sdQnD8Up5/sELvcvWQdd2u2dACVed6KR+VsEWqaJYxD3a6qdkE9QHpJf2iyYLk
ctfb5gIRAY0QzPfb/+khhXvRFgAcc5svUPFqCfVdLGzKy+t593Zbn72YAk8pknBH
ixDs8pRMwXwP0SgN1e8wUWobCWca9clHPyXPYcVfB1xQWBtzJaWj1g9TyZ3KxGFF
EVxX4LDIBGbcgFLdGEqgca2q1KVIUQ9kOpurw9nmUiJmnRczbE+DNtI1MNvcd+DN
0YHQLVK4OEttYLJjI8xalAaj1p5IDjX088qutZERN2I+26c018dM5wyyS/MoLxmF
HY+Iz82Zg69dik8C1euZOyFh7e6p40Cqd2IpuVuf09F0BGXTJsX2C/Ggrf1aK/KF
/rHelsOP/WJPrwFXFv8/nz9HLR9w2x1WX56Uo7oV6DHxsOXqiTzTNf/27sWBC9Vq
K2sf8znmoYMVhjuRnfCa0nwpWg/jRUVDDDEVXh1MNXPqp5Sk+vy+iXa1aHFZo3wr
JmJntxuxuyPfhRzai2CwiITqQVSUNnDMcB47jYrUS0wMstKH1Y+NGr81n9oRG53o
sW03pm4bQB+RfNqEGL0Z0pNcfcjBm/uqqhqJ3Ef0rTrsTGvfv+AKOdL4Ga1eTFRz
xscLsjpwq7RSv8wGDdD4GAlR1qaP0NOSj37uxNUaqHnnUTf0q8p87HqYR4cMvoci
Rqn7LUYri1aCRU65/9IpMhegVZKv7dpgkjow9J9vox02L4KTVb9w2w0b7sE6gJCt
Mbduieglz0ztczwtk0YzI+M31/LFiYFN5OgBgo5y4UomvTgZnfclseFdotQ/Y1uR
nRCbUVJ8qoOy//lTvSTz+ggwto42CHIcRVrl93wI2qTiYjo+wvgrq8cWs6IZtn4s
jZQeexelXXfEhddy041ugVONyU+s+kY23F3L5CNIcPQNZ9Tyox/mpQROKb4cDnNh
i2xaexxfAbUa9JJGGl0Bdeln50OSNwDxVqQVOPPQYLSCYutfV0JLNcHMDqiehwhj
38If6jl2v1zjhTU0tUUiFz+k+BEbOJgePydAIa8g0269vCdsxh3/LUbOKb0m6q8L
iB1ZSeXDX/iC4A0mO+rXvuQu2qI/BoXVRBbLIYmMjQYFE6JhNfsd0Oq0SVwdSQY9
55rLnK7UVhXH2IzBclRC33bVIZ/WHNpY1l3JhVqlwDYChVOIrr/4d5Szh4uSj4PO
A2XmQYePXdpXlF1ixiYbAHiZMNe7ndGNnYTxQuLJuKKaTexIK3uZUhW+54Yrre0a
qnIyBVcmVaM/M0vOrAm22zPnow6JW0ivjCsftz7A4dRRpr9AC6rgpyWUUYPJYuf4
w+HiKRzHaqn9tvChq8jMjJgaqDoba7sa0WG4gfXmHQsfN/bke1tZu4AMx9IE2LJF
aZe/7Id8+m7CgXGrkvHHphGeT0HAB9CHIcuYJzdgNBwyVGSazabWaeHwWpVCGwqZ
/EGavQ/ZbQA9NzoVq6aWKJh+Q5ep5HxjAhHCZDnHiD8JzPIUhDnoZUUYE5sfEb12
+ZdKBSyAkKv62QyGgn5IZssHco8F+XTkt9cCk8MkE7+6/bmfv2kVE99qAEBOm2rX
vEy1dHXhpdSCTVVXxYw/PB2syXoYfo2fxUwje2sfrScDkOezd03AkpFINMk83xFv
Jfb0t0uD0iqHp0Q/staWmOlX40Wg9IgROIx1HgKryaLN8vy6NGOhXHX2VlA4Arl9
GX2m21y3xHekRc5dG3PSONVPF++efQLwys/BHOFmI5X1Dln7BWpv/c5OHfI74R8h
tAuK9pd/ooApOsXrW+L3v2Th/H4bz6XD1xxoYsBiby2ncp/a4pFN0o0Okx2Ryn8i
l8qb9oOMAiEbiicRQTOg/kK5KL9IWtUYnY1sIX6BLaQZpDWugg1M2SFaqdhTXQ2n
XQosBiNXzpe3UauYqzjSPRbwOvHQgJZIbd0xWGE7fos+KPsKg+T4k5WIFrhZZpu5
S+cvZ+U3RZBwjzGrY9RLuqQoXppZL4cyW2MLwbPfqb7M+0rqE819gZ2fYNyHsUV2
fHj0cIO+FXMKxrYL1+9jFoqwyappwbuY2tmmhLQJKU+ZUplH4w0P7cDa20wWWio8
w+rVOAZaFIjD0hQMitYgEWQk3U5lgMP3JBT28IxkjAEN4XrqtyxFyGGI6fibdjU5
tH3QBvEOlieNpx/MkFO9ijsPR5LRHZu8qf96ksa8ItfLyncGJpgrpXpgs/S8yLUe
UgelAq4ZXB/IJta7WDYFg1aUul4Yu9GZ5amV01UKvSkAHU8RpAz9vS280DeEvxBB
kDUD60tsRK0L62jQ3/m6Vn70R1d+RENoMBarhI+mXBlKV+mfuAxHsJINASUhVbrz
00a+WnGiBxEIK6bxRFsFmotYjlOnEQHOMO/QUj1IUxdiMeWLue9XNPAhSfNmFh5n
TWsRvEibFsAv0xuAt9VSn9Eonc5g1iKEGJstoszENfHcqxpvDqXVna5Kj4W13U3N
IgXTOQ1FpTJ2x9/YAwPWQpuMgamqorAdempGnWJ/jUE0FIoZfna0D62jjZcy0Rx4
J4NDDxE87uVFwVs5hvYlqq3emswsx5qq2xSRU3Xk1rDNV2kEYO3Lo1ZPMQKezx4W
LyzY2mKwnxTppNnzPfQB3hDBGqL7wrz1N1IdUWSlZT713BL1gnddwa4Tv5qN0D60
yBAsBx+EBA7jzKfoQ5wWMwiKtGLfPU2XAzrBmXVN0tF1Qs89IwGP8OYX4//h6BRf
fT2za+TMBY4e6qZqYKCf1Wvwljq/gJRiXqef9rljbOV865MQ6jxLZ4bnIgy8vTMp
5Yfq3yIzL3zsS8speix6PK4gKVNAtSAC8VC8H0l1qZns5Pp2OGRul/8H2Hjy8IFj
61vVuT7GWuljjb4Srbu0FBze4Ug8tqdDxXQitZLvj51Oy2fXzQyDwUcpbDsPv5aE
bb4ndJ9LXxvThsVEavS7Ea0JFQuSScOzfU4RtvKwE1SmMUM2B3aSuRwQuzqJ7Yv9
GSg6fc9gZ01Pywm4Pc257z1ImAKigScWK4d8DFVGaUGDofF5wGaeGpdVh+92+lkC
Ta/W8wjOV69ytv2R4+gCFqHca+cKTU/k7y5lJS/v1Tunb/S6IiuOlRJ2y++adtBR
Ze2u9tLGsWJ3L4KjNyKbgdG4n0COA6fmnyUL1zCnBXZzH25Uvfm0CwAfnrvFNTfX
8gr8Qec9Ax/YCcs2g1bAoZLtHIHiE1P9BqYe8Jb8Y0IWjgZVO33yfcvqc2s1/FEc
2H9m0VJ+gPZ6TbMmHTso6EPiX59uoI5ahpji3/kK/fblkCk7CNY6Md7EsvCMZ1er
T+KPjsBhw0Npu7ZGpn5o5smLfqRZGXF8koIfSfoSF+mmnayMAjqXyu+I8WSN7gs5
M6AsBgaLaXn2lOye7p6t8urX1Tt4BGn1l3HLJTsay9AkHoqKSelAA9jxyaFh2Sip
ko/LAtUhwiUQ3l4+ooSuihyCZlcVRc1AMkPQ7k0jaDQOK/VamOgObcdOK4yj01r8
62CXqUfFHooCxK4VUsvy1sQVj6TjGxXvc2SlgMimxMAHFNg6zSztVaqDGPRe49op
7wCuW+lCHdUCTE7nLnObbIvOqh2DCAEXM/ZCYf6zXTjMUefVH/tB4hNvfFUQPeO4
s+fFpp7YaIJqUIPyNHcJrYJS7MkPUPF6V0g+tkTx/Ym+p0UMYKRCi4NjICr+sVIZ
WTUvU3KXtULYDLt/h62Y/E0mqfaUf6kC8X/H17CPl8MxiGwrV/4obrSGGlwSgAuc
EljZUh9fBMh5bfw+SHE1UnFsSAGYoVusOykUMfDeCZbBL08eQ/XMtpWko4++M4QC
cXn5M5RDqi4ExntZnLc5bdX0tVEPlcwie513sm48vOm/8FjZRLkjykSc4vvy1tjp
8f/B4vG2Hcqbw6UGwelVCCKkZTBrb/bJ5utl8A118Oinh/xocLzTDe8ZHuPAJBpi
gZsh9SKPU6kJUD4Jxi/lbkKph8oT0Dk7H+bPyqbR/uj3qN7pK2pcJNs41igk12LJ
0yrwp/0zVjPefaPgYjh9jvGAxjPGLcB826otRK3YZoBU+eZd1ZXes07HEHvTs19e
dNmTYcSSMeG30fZ9Z/nbHogbPZKTI/FRq9fFHiqfNZnFrKUp3RVrGU1HE9PutEmy
3Q3Y/x+mZ5vaCG4z8sW3R3ClVS6TtlP+mV5FwC121/rquILZqzPFI2Qorq8sJ19t
JNM6Zab3iBMNOpxoGan+XE0GyP5O6a7DktMbTwtRAvpZyZB80kCSfwNhxOrRHQPJ
uXOkJqfCKtpV7RO8GZPKJAxAeC2Z818m73LE1FOCiexCgJCMjkFgdRIAbSx6bb80
m78qidcrpjxbEtkyNBi/jNqgUCCL1utEw6YHEYkNd0TarzhE8JDvdY7p/Yc0IilH
/3dmq8nN/bsT5/N6a/ap/vNW5DCg1eBuY5a11Q61ptXQ+1PMU/1Luz/fMnT8KEj4
oBmhlRUggyfQJjjBGJuuebCHUTGCrEoZilcmqg/6IgWiKaAudUs8JRFGz+vRbRrq
nJtlz3U6ldcGrhz8y7vdC3Jt/xKZGts+vPr2okdImlOrXQK8SpD/jYH50Ham0wlm
b578PhqElwUwRPC2Y2sxE0nkqszYXzKIwszfNb3UR2RUkyTbMXG88kADlL6ssC06
0qtlGmSA20H21dCHmhFYfMp36+h6A6VUSo8OQ8cDkcX7GNdBNSeyqGcliD+DNbgl
+0GyWgyYV2c0Ndxo16dnP9IlVNM5oqagdb09DYLoVZPaSeDRFp+Llghtx5OM4t0d
4e3LznnZIgLI39x7baCaYxLk1M0UHMgj5F+cKLPgwgBUpQokALEl4JvSbaoG2etp
pGUHJY6xAYT5q3qgcgZ1yOH8nlJrutiPqEaZ0oi0EjoBFwkzq/gKYYaOeaOdcJS7
TcrwN5lBoWYxWB8ggyqq58vKP2KYFem+bofKdEF0eJUaOT/MOCdLd37qNjs/Fgpz
Pa8EK9wsgRkHQL6vv9TulEOyaDGlToWOVKnXTh3vtq4cw5HeXWRXDc5sU4JH1SBR
Tk+BEPQk1AbEGLtitJmIYv37DZ9MIiLDr+UMK+WgMgaulW/mxOVtpF1SAzUaLOtN
SLrC3wKUxv2/AtoWpoFk+8yRIhq+pbYRNAc4eHLgdlvdzJKjyxpwHnUaEBG2BAPM
hAPWFrhpT2AloSD2eaTXS6UfcDrnY3S0MwIqs2fEVBZClREo4yYtSGgmtH6EOmXF
uKSUW6oFNk/jMsYHbN2YRqrJN9H9HJZGAes16miyyXCza2eVgwKIj/OfTa5ANJ3U
6xcIVFRgxr/VGbBEi8pGZi1ora/LZN92GsyYXQ8Vt1Dqm1/PqNta1daS7g2opxNL
X2LQ57tpx4Qj2SbJgUULaMKwrdnvZG8tQWEooDJS+GP6P1r/07PRFXcBPivnXU9U
lDzOWMUvKnHL0kjHJ/LJXQteUr3opx8Ofm3saSRM+Ke/1YvewwB3pG0Hj/y2EjqN
PSuc7SnlWy/sYfoIU0CuUtZLrKtkQ29p1ssPpLOSNtjpwo+SE3oP9owEJQKBgXyi
EZ/osuejaHWtomfXR9MC93FQE9tTquCVru49u50TH8yadWDz/9RmaHUs1847rmOo
9unb1WU5SisPqCbbuhH4F78+quNK5zIytf3lLRzNygbjuJSyCJirQEWeVXw9r3UT
2Jhyy/1t/OxT9CNLjs2a3a9ANR4Rna6DoLh/LISZyWuij0QpLr1x3RKcXUA/wt1F
Pozp8+cNcgI7LlRVf+P7oDRY/3hagfQcKWoxszlxOFVPXtp5Io66fDkF53NVJEgH
+8UOOhjvASPdsKF3D7thDi7D2nrrMcZ3aMOOBOKMDch/iSJAvXaFBwBnC6OqsbUZ
lq5kV6mS/6vmm41FReXAl+m+7YOF0E57DyVzrGg0M4Er1FMuNPa4zRJD2pu7nAHR
4pepFY5ygNj/sKABFygr6hEHRnvDXAJQI/CBD0tmJIxH/whbfNCuUp19IGOPELUd
bZaS0H1AN4/vbUm1lkpj9BiNXhz8uGJM7RVwbbS9z30Xl68JkJsivxYmCXlNj/ty
pHuVaRoyAZChT9s83tEajNBDj/VkIRp7Eg9SlHXJiGpcTLaByWBHjUKgx8vQHPLu
LKvHPt64gyI4x79Kqc3BP/YSi8gRVffV9mDAuB+pNQgYR2WPkKrImdu6Ru5yV+MP
W0AkjqxhM7l6G7S4nVd3xhYIHAZJpfR5L9fsoYzvKXJVoZq8EZMuqSuj4AJlmhfy
Nal7t4AvTscZvfkwACR7gDDuFDRnb265oK6uoUacMimnKk4Lsr+DwycHXSwW5Skj
Kd+EIFoVVFsEWH+v8pbEe1u4r3NnpB74ybHaRRFpxKxSeEQZQTFxt1rVk574coVA
+e5UewMJ2m7noBYa1BVY+J6i18elC4tQ85RiUc7J3T3xif+RQgT/YSOGtPIqmxjj
pxTIf5nc6i5+ghRD/A7xPoE0zP3X3M/ClmWr8ccG88nuIjDUm0ZhnzthWmtdnnvo
BJH5HfP19BrTAS1mdm6clpoPCYcyeaT9Wlc/wGsd+0rtRLGChySDr0rEp76DLfPj
5pAjoJ8JEM02tNaE9zP04cy5TXHnqIhXuVzfmrB/5hxfYO3Zo4vvUH2UoTnvde8p
6gE3DIDiqE8Zo6XQjYcrs9bXKcqOEdjqiU0wEjCUO5/STvbOsueDER8z6SNaI8TG
7s1CnNEN8M4xtOKdQzHFxPm9NbRAJ/2Z2MF8cvMoF3iCPOly6d3M5Umu0dKSd2a/
fYVg8H+rxNsVGcAyMVoAqo0mS4qvKBYcWXhpyMoLYy/tEDLJmcg+fQzHFkDaXTUc
cwQ/Bdz2+RjxVrD1fPOe8s6XqqEATxtSPa+HxiKCXWC9XeQG+7Sf4dMXuGwlS63q
xHcnrMP0wevoNYGfDpEzqgE07Qp0bcb3OeNnc291ClFSScBxbIqF5UBOLY2DKQrp
nxqGWN9CzHN5ycoYAuoVac0QDa40oOibNlfJUT3GmfW6GZ3eIv7fCrqDPiQUYbLg
9M1Z9sDIeXzsWBmvF6fUTIe6WjwJPjD0ONQtp65O92Q6q+u9aerbPTVD/+Gm0Q2U
NWurcIDwsjvKKzf9L+P+j+Bvvh6ho0wThSBvi0jhaXQdOA77ebxOUy9has4tdXku
jHRDJPnOW5+VuTqgEnTW4uULN25RRa3l3yZUVVdpH9ndsnDZ2NUDBc4Y5nqoaToY
46JKOLvyAG6HhGqhgxhToJLgbrqrh0ZlFIzQxym32Hpf2fWEqoq1AvI0IoGGbDgL
8E3m/3XVPDQY4b55q7DO1rAR+ZY3yDjnUCB3f6+3nZue0F3kfwy9Cz/XSiPHo1n0
+HW4Hq/PyTPr+eXcbFYv46xDCZFLx7NxHKiSM5RY9fQonUcsw7tMXhuyhR+g/kY2
5Hb4diRW771C1wdPf4jpqSpGSA21axyuoP/SjNfbr8XHGa9838vDRmRPRl+JN0XS
ARc0NHv0k3YR70INntHGu24czQC8O6b0K6YujC4npJC+DPzulSPC5ZDQ3qheBHXm
lXFykMUWAkUObqyKJDb6vPeg55pJO71tXT+nVXdEn5N/RMaX6XKNZnqtDPsUAkBI
3ay4/tpfbx3G9yVFkwys8fMbSggD9l2I2ZMX88QyeHuSdNM2TgXguL2MMIt1b9eB
xPenIDduHuCtfqIuX/J6KU1vLs5BQi/edS7wzLVaJ6kywKoLt61shJtS7oOB4A7r
5+TCcHiFFiLVI6Yf+AD3Po5rcMG6wlMnhw9mOKBQmritKM3sK8jPAEI08Xhrwrsa
Hlkxjpqx7lhlbVLJiG6G32APyXAZs4e8lXLzfcjW5NeUvbUc0wVPSnYizWR5HjSS
fsAcpPcgazE+M4dHjQI11E73WURH3QErtuFLIQG0my6VrbdOhcc5pcPTqrWF8oKj
gPX3uAKc6r5ngp4LACh/+aMbhDaUpy/7E+VA44wFE1BvkUD2N3suJgt+qbGF1e/5
Vcm69Hy0eonW+OGJgnKLqyqwVcxAVs7KzH0pVk+MQ2wDUwDqvoNc28cTOYQoXnle
qZF5LhMAPhlmIHrpLV8BNHbttZ+j/Yli7syLyhUSu/xYNdN+8XbTPx4FQDp51TH1
MhGlLiosQ9U5HKhY4qKH2xfn1YUQnOIE88sH8TnH7WZkDetd9uZQurI6w36ifTGg
hTpRvb/8O8WCTEQ+Ss0AeEzfmXoJXMcCOrOXqIOshGWR429ddz3oZdMlX5iSUl0q
7tAmyIGG7FFxXln12PxSuezlQ+qiGu6UE6PX464vK9qz7WEV8b41IXLtHKb6EjTw
W8bWR7TQcrLoAapv5GdeD+1+L0gSbfrw1V5K0sqXdduo7TXiOM6LAS9hOXHfpnkB
wA546Aezo6vs877bQDlSMurP47y0DaGkSbjZR3P33H8CU9oJxlcf+OxjABCx1zdH
oqxD37vOGgmEo5Auxqmpgyz+pi5rMdzO4pE5VtuGsoPQBl5l89/a2g4QXZ2VzZH7
TNbGQgg6MEOVAsaufW2TpRY93Ta/D0QoJDVU3kApGTBOOadj9g+m0XoGBAPIPxMU
t8Gxf+44fKAh3Ur65v9E8yQbs6vQ5hr4yor7Jdwn4GYqRcHBuWK6kcNSU2/vCWL3
I9OnFF+spwSkT2YBEk/xpTxSZ1hsnoziMqJSTPVXEwLjSiE7VYnstK90vr0DJBEi
CYKOIXmbeg0lypVhMKYKQnq8ZsvKIAe+Jp8LFpcCiNbRlaUI8UDK0OG2tadOIOan
/TNZejOxNRHe1Lq9ySZnipKipqsQAak3ZA9RzZEcSN2UdYTJ3j46CvvKQg4tHn8U
ty0t/0WjHUA6xrEUTUB+XrxgKpcOmdEdLOt9rIotejaw+HdghLtUfm/onClGrKtN
18hvgdI/VPajIfdMtAy6VNm/Xb7bmgAuGvIJsMUptf/kP6L6ibEihMShxRBTfAEb
y0Gg7SzvjQBjpHjebMCmvr2rx3C7A1vA7/zr/xFlBxBO7wPKHJoJjy1xgfCPZJa9
TqvKFKAnxYFeLL4C7iZaGxcP7auJyZ0Bs8Qxm83Udcx/oXtDuVMOa0Fg2eH5elgg
PYxzjznO0Qb3okudDr/qoxhQGYjoauRUOcIp3Tz8JJPG4S4oHtxpHJ7RKxiYbd9R
1LD4qf27EjSsM/CZolSlF3Y7zopBVcJAhtZkEfIexhBvMrTp7e7AQTpl1TYpB0J1
ieBMOJtrIL2vuPEWKpBeFhldZEu4pyrdXQElmpuMuGc0ypkbsYy04zAV56sUlBC/
7IaRsy7VUv62RDMyJbozD1KaXhSYuGWfUaFAxoNajil8IhsOSy+Ljs0iw6HRgayH
COsw2q8cLYRF5mdX5KYOSblMq6QLEOm2fQW1s2i6jGEomjUDmJgQ59bm0A7uJZ5P
XGONSRBlKxliXTgK2r2D8Nij9Y2v7l0RQ0gYkN1RMEyYZ4U4QCfY3tOK68vdhhD/
Gfy2+lDeP3HnYMv/e4eDvhUfhZKxnCzIFQAvJ0t7FJJbKO0KdfVof8xMySKvDx3B
jaKk7vFyCBy54McaU33PPhGRrBQ8wq0gphTwd/j5vS3aOmQJP08g09QhblFhQJTc
9RAxAEgnba4z+g11Pd7weFtOmWZDOfRZ23NvOyrvY+ImHPLsPLZw7xPzJKgEjIao
nIazhQbQ+nLPVg/cGxsPC9BBoDVI20Hf/eEy56p+tklpTIufzd+1jRgKwXEZeyuX
xs0iGoUDUFf62lavsRWgw5LE9+c2fx8S35YEaeZqHIsRMQuUumnfusR/OwwlO3bm
9CpINfjJhiv2boIEB5YkkLSoYB81ZaUJ9e1puV+F51hqzW6qry+e8GROls5jlsZb
GE18+s9cyLwFGwkPtb2hpER/XSUG1N178GvmUkPXoMYqhYXF6XuYuu7lJB+g39LJ
7JdIw0ivx1ZSdFitbHV9FqMrgW9CcNw/xpy5q10e1vs7CiFnzAGloLfV5jrUFa0p
+7FqHEdJjRwYGrHyuyZMC7UldxiqfxRkXsky6/wy7vaBcxkalxqDOfKnaZ0OESPp
mIosDRkKm09+7afajp/R752w2aZbynXLonyOTGQuIzEY99x+ScuuoH+oHbwV9fJP
fXpwQSq5gI9Boaf8PONXBVA/cLEY488yXeP2+DBAv6cp6nfWDJmqP9rOus9AA0ds
Y0ML+XNRVQFmJgMbphbcx9w4nm+yAIgkpfsy7e1VCjNCTeK6zLZa9HJ5TC0hBR2G
76rXk5nCBLqRO2WrPqkW0wdbalZgtegkvF/XgwvkIL70j4WcYcOJmsXAayGX4AF6
yjthHu/E5c5wwW8gRQ3f8+rHvE+3PnELzFS774c9fjx2C7rCKQv5eSEu4o2XJ33u
2MCMq4v4x/NyWxWkJfXpWB0H3hl2auWhpV3l9i/bcaUfD6VW18TzvJtMjjeLECw6
6rpmqYQmTV0Qvg0tmWll1c9Xmjy16xHFqw+y5iCfMjpV7RliE6OgTFXyv5BgRYfr
M+G/nNxirnCDFiInYA3FrtsGcPvOYCoJVq9mq+zO3fqhO81HESzo8Z7ayFXBz49N
WIFsn3RQ9EcAL0iwSp6Gzbd2B3iv3Mq9U8JhnfGOGTk3Omm0oC9fcE6QrFc3/HKE
vbJEcqlz6Rxp5lCE9Ul/Ky2MaqqyoN31zwUtRBj4rsknl1sA94RFA1UmK+ude/Rx
g5JXsx/SqOmBOaRnQsFugUCwBWBaMfnhXHlGig5xcUQ68l5AhjD/FT+r0J3dJcAY
WS+BC8PzGRoZsUdF1GYu5DD0hMyI51d3gn3cCn+4/2mntyIywok8XEklExexEYrT
AhLODxCnQB+DtWILFj2m9Xyv/Esml56RJm5WTsfyRWZx1Ks+10nMkB4pMEc2y74I
rRDBwvf1ZrOB/t7obBG4Peuhno9xxT3Z3fpAek0oEDvsCRJvU6DXjZlUEqF+QQrW
dbQHg0zPgZvScY+BBigmqeU6u+yJcNT0wpKmbXSW2jRZ1QhbkhAuq8tQqCN1Pbzu
LDYsJ31V3cdxeWHr/aUW8i++KiIO42xzxPd/RV73323+Tdo8O7aj6qj2V2EQXY6w
dYNArVKTXsxDAdo1eVFyUBi6NGD7SCBU6CshimqjQa496uzh6VvsG/DCP8klgCoq
xmM/YBX6TWyssfVAdeRap3B1M8fG93ojbVRATthI8IbDP9bRY44Q9DSnS8JgnALI
QHeuy3fNC/o0Kr/ca26WjRZiI7mmmWY4Ta0IgsUraalaFPJGM4T2kXM/Dg+xksQR
wE0k5e5x8wXZuji3aj9BouzcHEPPF88JlEEMMTVZ05xYltmOBQmoAN6s5ewk1uKo
VUUIcDgbiIqcoBnFFSS16B1n4Feriv8J7fDBP/x9lBL5Y0+2wESF/tyHh7YTOn/l
60MI4DDwphejEv5Lo5U8E2UEnJhyzlfTg4aev9ZdGxoj4Mabigpkf6CriSfu9bMG
uph1jYIFvKASunoUDHcpNXeZ11nUCkq94snXsGPpr/1ZbI4Vf0nSGp78tuRzTFDO
PgVyayBXtiRnWK1/xDDdWTGLWOv4jjVdDehtwoXAH2tEN/9GVSCZ6SVOJT5jQf25
ajpv72AMtI+YUjshMS8NRVVQbeN5+wvqX3Q98hiN9WHkqTfYznjWhxy7rw9hs09I
DfEGAiUNBkE9SjG4VyuQ7onXFMES8lSdlHs2JXgDg+q6ObDnh6evYgvthQeos3p0
JRrmECUBy95agLCWe1Dkk3pGRbrlKaYa8lEZkEcU5exYMfcdkucaMY+PBhOgYt1u
/jFWA35Hh2XmXbaK/AVoYeGSBQrZ+jann9M8i00quCrWDQjE98RyGEMEuZ5TZGJK
iPMFHHbfCZnYDHqn3UOeZJzxrcB1t5O9FMAodiRIkUherjPO6kCqdXCrHZPmYkCg
iWNeVme8uhnNYo2Mvfaor3suCPKGdIp+w+1+tg8d00QrPCAu5/rHFrfOESyT4h+o
MknS7jeE3R80x5uC1vNPGScvrlWlnxEIQDbt/sag6TiT7OYkCSUNCN7Gg1KLmfiF
4V2zWnmYIZTTZFwQZ8QrofrZqIJlslroJL9d9Q36rikxbv9shCvNxgzExXLs6nE2
QURnOxPNFsUpw8y+eOfuxXXXMK3zwMUTqqo6dgbjihJnXQlGBfiFEOelFlwStRwE
h2whAOXOYuYeeROC68ucihtlz5pXEgNhwiwKHHOXM0bmIYGQE8RF272dMPOQYuCn
etdFMr1YVvrUSk70riuzGdT1W+bAkh5LIWVkOWurhG4p/dS85BnfL2YVPwtenQbf
FKth/XiRwSxro5ZIyFiTyXH+9BD2hJNCwdX1nLbH1G4HqXGDoFrMOwn5WeykpbxA
E92Z1udYP0FJOhQXQrQUktd2v2QlHZUOA1SUjF0YUnqhnsKBVL0hWsGBNgG1YVvv
yINY+thQWc10j3u3OTdXlqj3enZe9+WDHuhUAQdwsJrYgIinuRoYi5nSsLEJbUfY
HAkV1zrrvxsH+247UoDgi0OwLMFZZWigQBIV6TYg3ZXC2F6/zSrqjv20R4XIsFwX
Dyojttow4hm5JCNuejdUfqZkhGgwGZo8AMW34zQO6wXmRM2sGItud8ZP8B4CdC5Q
QKxYgCjBq/udtxuY7FDYgl4vvo01iU1PxC912F8XIAHo2AOYzjBR3D3xzylg8WZY
9iRtNOKOK1SitOJkhbTf24k5g+JtPqN3PemjpUQN5x6Oopm+/OV8B4jfXxZ3apWl
odRFbBk2LEtcyDELQoSgXj3J3MadRWSSAmmSeTJ/n7ibQaOASC7G2K/IkAa2S3Sc
mxy8vkWfVgMU9TCkEx8+mJMmrDAvnYEjYybioOGZippOPh5YsOMzYltphE2KZ8OF
P/loo1/Ou8NR4kDbuxRp1Si/vpYS5t68tANngOlI97xJMQ5hL90/t4uGiMtZzt83
Q1b5fNss96La+XAk5IpBkZf+EvJw4Orp5spP3oAv+/85x9yurbWFddelFyy5YNxp
J5hyyiHTgBSckKgMdiduo+0m9W9rUvJis/StFEshrqWZ4ltc0F9ld2JcO8JrkAoY
ohtq5PkwxyaNBmPcCIMRUkiXfqZQpR/1bLCuR9eLAjcMneAvCAwRSJqCxZAW0Qio
rEnQvXA6ZXw3GgcCbhOoH+FRzSw2LkPJW15ut7aKWSXOppi0TYLI3ClekQDYtQQj
yuIKQKE9Lusy8zFb0pPHSAub1DEXAa1YrbJEiqb6ck+4yfv6hIeCLfD3Ww9V0FWC
QHPen7w/OY/PpwImYzsoe5qm+Mg3+Tk0pARmzM/nILbZnSD0VFHdzTInv9gxN5rg
0g4lackcEkT703y0N4/dA06NSZnuhsOkGVnQ+5u5vVPb+MCOK/Gg9f6VrfuJtoQQ
K2TdjThOh09ewWxdwOmiPSZH383N4My2w2UeS/yUHEtGxWo0keiqlC9JcapIVGdw
8RLFdYcw/gV2r8r/zDSE+CHlcF8myjCxs70NVzK/VGKkheYtzOp0fjL7sCXS/g1g
A+sMEjJBKXr/KYtdtduljIqwEC4jCa2wOEbSTCiKJyitrv9lSs7sZVf13Hey4IH5
bIEO4RF/iesOGy2fN2dCrLgpCQ44LkbUUqd2lk0PYQIlZbctpZwH5BqdxlvlJlBU
lvxt+kXKN3ypci64L1qYcC1ELCBZADaqzjjJk/dF0rfBJlQzjIX9eOhTcOa/MvoO
gyZ+FaDPT3H3TohA7iajc00saOtWTFvcEI/2ifLAa7v8HWyMLPupAUykxk6lZu4T
HaJNjgk5hBaO0Fp2hXeQ+TAC2vflEBvDG3TZV5QhC6MxDhqvNoE7PX0s4fO2ZK6j
mrtmX/rsisvJ7iQOOJbw/dwPoyEeP2rt8TBv6IjYoRAGV8Paga33vE/6oerNbp7/
D8HDEh7Y8+OtlbPYLd67KE7tDirJDjfaKB25r0l9TY8L/BMRqoRc87xI3On/CokX
2p8HfxfeqbCaFWNqPysgxofcdeWg2wqLIHPO9b+7ZmPQEdIV8AKwSx9VKJGu2IbU
cA/8sKzXpBovvo/K9xLyJdtMO3mKeN15it03HanVfMQWZ151SEH84IyhCU4mTIPs
y+hhMqMAfbteYYnVVJ9qi4shDxFWUBsN6w05Ng3JuceM2LRt69ns0ga4HF+nLGd/
J7s7pipZgfTt+yniWq28gsfmqjzAtqrVOHRr8wBKvyPqMzuOohKCtvESYYmrGM7Y
giKFn/iDU6FS2oC0ZWxugKsZIG+qsAc/Y9jVyBcR2EqeJ6Ek/xtB7f49P12CHo4X
AJRt0J9A6WwYXl1K24LQ442TrZ8mFs8zhZF8/vwvv/onf7c20PGRCXGpWwcdWvKN
kiRqcYDTQ1tAcINHSt1GuaQjQ1/FKOwwaCJKajQXCQGUGy7MgsTdKGtafOvz0Xor
jrXnrjVakT9sccoVVKpVY21i5c6Q7vOVDZDR5hgECMy2zLX35KqYLWuKD6n0fhU5
p/aX2T2s4D4fnX7szstfj0AgKZ5fQyeagobhU3ABWCOPTDiL69tMtlEmt/pTIteB
T723Evw7izqrgarPFZ/Y/nWNPIPxpw9wE8m+GiBC7q9Cf6RwdvsBQAMSEy9uunJz
EPIqqeKpg8ZNO5APd5JKsrm7Ig+KZ/K1MLoFdV+K7ISIf+WEiVu0MTI+juSb7vd6
XJ72zhFkNJSsJ6txPunYVgfYljo/pNfm9CaJ/LbASO8kRT7xw25uDVm1KPjJGBEW
fjBojEKBIZBsFs2xRBNjN4KWMfR1IJZG7Prdj06nBaV42JrzvFet6Yg6dSL+IbMd
PYi2vaZfPT8B5SlHHHkfSkLk8GAgUgj++ylGIRFK+PoDVFICe79BCECtUehO+hil
zf63nC1I9DTOniRpeQ1Ie8hPkaYvvfw3a+HaVcVMLOQ5xIl9kJJrh6dpUkhByMwN
KXiyu9x+a3wRvLpj1YgRahLWIbP5oERQycC1j9CjpAeaat6MLWj3n69Uo1CzRZEz
mnWdXqSGQOlY07YT+DfAt3yh/FQ5xRPEg8d2CjKNZIQqf3Yo/0RPiFOOOmAEZ+Pg
ygtpwvAEipiHbQk12oRnWYR4zPGJuxspouCI0G1SaUle0btlMINZu9orqjn2WpQg
Mj/KpApwu3Nz3yo0yZlQrFB9zyp2PihHSyDDkPXgrRBPKlXriwfwNHhKoO8GQ5au
JzGTsdNoydult8JwcgAxybMVTSiRBKYflFltu0OsPUPmfAJdJZyHUTY0FTdKrdPS
rCKptEp7OpSG5fT4wVIK2XUgABn3I35WKaJPy5Rb+RLWDkDKOUfsRBbzrH6337ux
x528UDJIurHDRp2D7Sur64gtraXc5qm1vXv9PIr4Zt+Loi18++hCiOztba+nI7GO
s+eRoX5VDfjv2QIWHZFO86h6435gGT6xBOiQXLjraL1K1aOKBq2gNEcop7wTbrs7
XmE3BXjC3wUttY6wUGdZw7qPU1b8ClgSDB9pOz+jefQL1PPPG03fPh1UGSoOJdMD
XZ68t1LkGVVQ2qGBiDGvahGWwipcv6HtFNRrmh/AmaNytCY00Mqp2Zjy0Y/Slc0D
X8B4QfMmSxQ7h+OCh8X36IkaYw0O15SRu7ZIc87WReifcSUTIGkkCA/BxENw282L
pejrs5DyKJJKv9hYnko8Bnbt2K+UqYxeJzvFq9jZntz+4nXZ1mOE7SxQ1aUB87xe
kksSt1tKmLRE5G0M8VrNDVmJ3hm/bUF0NYwTtErdI1Naya8p9Z+C4QK4sOfZnqfn
oEUnpiet8qMQpabvR8eLjVxupNglEnoEm4m9HV7+aSY/a2zpGb9aYA0kpwjMXacv
te2CnH7gnUNV/9fzLRmoHZIuaOWew2AwKuAXjfpKhR5N1gxNXKJAUUWWHD4GHulR
7UOsOzsue+dIH/B6HhRBIO9sg5zIDm581yPj8k2xDZFqQsrwZR8VS0chmwnRcmDL
klv6TX8lXS+9bO6zHAG0t0TktH2q6R69BG/i4OW1qwwMOk5yPgtMWep+Tr3psfGo
sH6QC/kesUchePcPgmz2FQmxGffjyBjN0cMoXzdrYD8+Vk2YMP4UkzzyH1xAYX99
BOgdnFaRbnaFT/mkk162ZoQMFEo3CfICzV4/egcshFxfe0EqoolL8wqQYnMEdzHz
XJbM915DJ5C/hcviEl/ZZvwm+r0mtziGxk7oew0sHrwM7Wri8asNkwuXUVsKIKJF
PwvXT0/1+R9GVuPTWM4A4+/P+qlGVPN70RS1FfL1vaG5mSgXS7y/W3bb5Qsf71OX
iU2MpLt66qzIjbgPYCsgEEHUqZaK9Vh1i95zxlWVSd7SfsXv4AaDuVRNPUnErgA7
rvstSYyPpWUKfb3ngBT7DfLLuPG2DUTnxsghd3bJLxzoSZCpLNqJFROcK7c8iAWF
PyUXyFCmHJVexTMeWQJ7fuC5tTdMXmX5yIzXhPKbvMcnTjWr+j/RkqnvzXesZH+F
xMEFlQr6ML+kIVeEvnkITUE8jI01TyPrYmGjT172SYRUAU+vtFMNyDt9djrOzlSj
mDoWD6U6FO8hDyQNMIrkTUyo1ltsAoHz+J4g5OWWmfv3lhdwdCPnZB+icbLHblq6
vxJZCYiPRe6oZzqUfM29bVjGfqBQafuIavTe3lVhdLnMBIEcfWy1ZidE0XSRGKoT
nj5ncQpXBdkUYjy7JfNMX91eiJiOwxULOOJtMFFeWD5o+isKiuowgtz2YomcSuek
Ew2EPqCCCnaaF6nbuMHz+q2GUFTWXn7g4CtBp5A1xgwICF2HqiLVn2eikRFRcHjs
p3eYDnyxsZvTXyoP5dobnY3/c35TJSP19uVtudYPONHVMjE8nbVkBYt8bqWN9Vsh
eKzhyaO1AttXdDg3p1btujvxHfW2IeQ7ZrleznxSGeeOzw5c+Y6/YhEyMqWzEbAD
XTEcJVtJ+CniSLhx52f2N/dFuonBeHfgF5tJ52USQhZ9m4gLANoCY4LdZIiUelHg
P9Xl9i0QVr5//HhOo+JXPhdUiKDnApD2+1SYqEXAJdfwrr/JzrZNwYRqDA9j0XVe
ZEB9Lk45Kqcyjvdnbaaly9FDRn15Euqb/rrnLp79pY46IbAdeLPPGEB3k/nUH3g0
9n4ktqjOUetNxS2+aFneDHrzuffHsDMGRBdXIDDGGKx5HhbdDo62VNmuUojE7GI8
6Gn8bCVYe/VHRI+KWVJdEusZHqF5QJp0/86UuKV8iS7aZDrt16JkeALJpvimSpBP
jOvLmhB0iRB5G9y14THx9w+CKmwwAW6bj3kr34jc6m/UFhh2+BGQ2Mh2QpEmKe8G
XjSSSznPvn/CxApWvhhL7WqYuBRlUf81A8CMhqCoov6foWUnL+wN5vd6i/v2Evk+
a89rAhaswftM401zI/DPVSyRdbmbhyy6kPHgDmazAlc9J6yqhxn+8ThWZDDwtX/k
TEKm/qBCSKKrHl8FAwDQR/h8tCBYiH8jlrm3zF2hT8LFiKuVmKymAvv3kGjpf7n9
UFPghpenNTL8VFpMY5N1YzGGMzyf0TFgK+kCfykmLjHLaltliJoc20iUemrQGr2i
altMfnt6D7soGudh4Wm8KNkkvPjqbR9VUvgywPz7h9f4pOaZxf+RyOMxFJbwCRgH
cUCVE6oP866FmUlPhw928nU/AqaP2idEEM7m3dTblmSDyXvNzdyVFIBmau7suML2
CN0HaXRzd5m233v8nJLZuCzQqhamUmyld69BKaPyLFO2AZ86lMr6xJ2Dh3/yISUg
MEvJrX48ZT3h3hK50SbDFeucYSoXkD+KfFFYkj++dzvLNwitaM6NR4VCWY3+sk8y
0Rn3kTmDb5W55muF2ydfCBBCH1FdsAn67F/66r/Rcxh0nH8/LYTm+STdiKom1NWO
wbidACEDeP7pozxAzBOZlIEir67ma7+4t3EFk4jQpoAfhxmfDk+MNw1SevkUjWcF
qtpAmUYsGm2GpbyU7e4esPoaK8o5frY/vmlEy7XdG0Vc0oKLWkCnt0FASmJzwd67
ZnoO1VrLRRn5u9wZW8gilu7hGitYyGeO1+eIVuJhwcLKFjdS2V95nCX7efupj45t
kzQysiSt/RlHpDNUdhm9XB5LSlbAtHZb3q6zANLPtsx3bR/xZCNfBD9bHbMFzXre
KXmt1iADWbbqUbXo3AG6OclDKGNXTgAzFdk4ft2dgGDweG03ZQ5K299PAzOhcWBa
fzJtqK7Rp17tEgL92YedO6fUMd0vl6++0EX84dW6y48KjqTDikG4pA9xDdvE69DL
CU94zuP+tR085mSfjG9fQ2kc1SjkPy2NfCIz+G6TfAHeYwTHxdGyRDdt2okkzQpu
2cpMAbnY6ZZqPmnDEtqO9mnzXcvLGh+2L6c0yn6S3E1xEdwqqFnOD2eBpxRuJJHZ
PbAn5QVuJebFLiupOqY2rIWQaGabSKMd0UX/FaNkOpTs8ySGCXRQ8adB06ffQ75H
YrpeXf/lRUz1DuFdQReA46yn1ilNNRckUHSPYktySKFuCN86+/+u6Q7fmL6MeYYF
CJ6sBpKC3fI2LpZ8RP1MQ2TBFQHoCU+RjtpwviuNpWYrTlRTNpUQH7HxdKfPn3SW
zA6nJjk6BCN/RAHhSSGHv1KFf3eLiaXP3PHSh5hSfiSyzDECHGUe/2fcLAPel2CU
pOrAttshSDEJYCdSYHODkFLUIBg7wPcDs6uebDwAf6h4zKs1p1dsoYxs4/JZ6ZXv
7ppqsFuuCOXI3wSOoQgsm6IMOk3dgVgVqly8aJdWcqKf4CWjliEtyppYF20H1IEB
Itk9AeXj5fxM8iKyDlotzB3V5D4aUlcMDnhnBuQIAlZRRrD0yz/k9CJpq+kd4P5M
YKkSZL4IzUQv1dc4NJE0S1u6+ve/YlToJ6m5Lo5qcDhJE+rO/zrkk+nzM91d2UVO
b1yNsYLZLnbtSHFUsimC5P2TvOpcTQ6WBWLWGd0dRQVZ7AeQvj3a0iZUf3QMBpBv
lwFCSZLEWpwxRT0c0fzMJCsQxAjb5nM+k2ta3yvra6zYrY/ximlr6qD4y3NuNNRB
iSq5qiGC2guSGX1RxkHNuRcaRSKV86tu3E305cDhUcaFmzDr67gUY5+/AFT50WjQ
kIAa+8eBqU7V7CPDOQdlof/fedOzP8pMEPFgycaIq5WWsJCmg1PXvF4H06dqpUXG
YeA7sqVNcYZA4Ol68CKGs8V9sjRmqUiRqD+IVhAoS1N/aQyDDgC/8Kc103o4OlyF
HGe/uKFA13mDFDojafnLxfEdWEim/ZRb+Ly0CR1sGDqiJJFmhF7vbq2kK5Fz+Dy7
3eTZ4v7I37e990gr+C6M1n5GE3eZICzOWg3I9wQ2250X55dcURtrIg1TftsxcXHx
hamR1ZgEJscFCq3OEs5j+zeRY+yf0jL02KSaSDvrYTNnPvn7+6osAwz+YBlOMcOm
qxHDiERKlksd8BX16dsWGp1GeNNaJxuhBhqfT+yg2w+2roYveB4qLA/66KLgPHvA
ft8ahQNorWPFwjEHBuzgmwkjY4CIhu5Eo17s//eWASuifXC7OWMbzr+weDVTSTYS
KWby9iYiJdMPoxve942Zt9SM4UcEQXq9wDOj+dsOmEiBfp9/hMUl7Kl9GK2vY/AR
e9IjKat+gLDsvsSFjNEgiU3F1BJvmqM2qEysb0qCeuZSD1i3EmM6rAfn5kHJbCaX
679/ehUUT3rdW+KkXw04OcJ/19MX8pb0yGK45Oj8+l3tIsupbgPQqpcbnqwRlLIG
P5vokWMHMIOeQh0XooxVpInY1NZtc94nYJGiOmYClEg0dtbTiDvFtj9dFY/tivVc
JpD1OJjz73MyuusdUNevPumunx2LkEyAfEkbQ3QYllP1tZRWLHoISSjDeIOwbJZ2
D1fAHTjPF7yga2o2VfG2xkA4uIHixcY8Ndss23UVfN3t0vTvOVDWKJigFmyAldDK
8pL09m3hb38ULoQwEvT2uFJ6I+SpvjHSPp6JwZQNiAmwFCYNjA9nKiuhbv8Hu3/i
C7QEHy+I6hOSPmW6hJX2HaxYTh88WjxDf5VcxZrLjrQ+D7NoD7s0ocpfzjgJOZGG
T9GNgsv2cp8QFJAGnmaBF4Lv835NXnbQqWM2o6V7Q1cy6ICvWFgdAPOT7lKifzY9
Ziv7kyPYO2fhpUMgx1eO9EHTfEUHg9gi58oRnOxMzGi91rJ09FJIpP6IBbzBu98+
ISSUpm1baKI4hMPJXXECNd1r6b64LdgoQTsGKc6k21w+VV3dGSbDDnioLFFVWZ+6
aIDp8ahcGQErJSvlZM6OicJ1++aLgiyPngAPNGNwYLY6xGNjA6gy44UU69cPLEkv
K9invMBSMHiBQQHzc7XuYqmDjc5WRZSnuPR8+m5oVvqQws6Lj/y8fvi41ppfwBe+
6lIJrSEW2V1Fn4m3VysgzktA6idumjWDGnrLl0+rAYdXN0mHD0OTQBkM+MkxgXHy
OPsqqe+BwqqmDynZXYVrBodioMCkd1u8T5OQkZzJd/7Jlc7r+aTfx9yEgKlHL88Q
lhe5Fiiu16HSl+RuUCAjDAsn59nag2bh+0s4lCtFrIOpN/LrzgoxrHz+8KQJyWf5
4BF3hvfRMGeioVHQzA+s2rWz9Gy8fiNCx6IBLND0gRHaEKtoD3YBptOI9deqYrqT
wyNtoblhTwKsFFuKLFIG95dT05eiNBYchL9i4lnqJuBReDUqPp1QXpYUNxDpjNpA
nBFFMb+JcJ3aJuF+xuWZEEzdyV7S6IH1fA4/iC3TiUdhBFKaJfFEhF60Ts8h9Mfq
YyyfJ+gIL3pk4Cs/pnwrc1ztDBZxhNQeK+DQY5nrshe5LTXcBLypuJ5axmaYcZBb
bQZfPHP8QlK7Fhy7urzl+fZ2o7orVim0CF9kJBJk+bnKKKxB0VxSZmobW8vScI9o
6YgPs3eJer8wmj41FlSmS51nNWAjVgUN1ENHIEKRCjQcCYz1Bty+wfAjRvtQZvnI
NWmZUUCNKOROf67oUlNE5F3f81qJRurNglKtdpcaO2C5chTkT3s2SKHlJoDr5MeQ
vKKeD3Gxbeg+jRr//1QhsH4b8Wy5e20rVM4gKyhC5+97diRpyV6aclx9aSN6K661
iEY5u4et684/SkRn8/4jc2t0/NYm+XSHHTgst9dB98WBa3J5P2riuTSKhICHK6tp
tNCKeDoTDOeR8LmsjPKTWyAFuamWxESKiIlcVzyZAXBZgEUoCVB+gN4pVQ16A7gy
YZF6/1jh9sHJ6+uVg2NpEhrH+TWD2J0PY8VrEn7d1eQjMyxkuuUi6NxUsrP60cea
ub2RrwAJpBIihmbg87o4Slo4pmafMPS5DsNT1UYXwRNXqS0mOsdYbHSu0KVIE8Mc
wn8JEaVlH3yK64F9fkCVKMZXu2ktz+ePW2FmBP18kU+E2s3LNfqCiYx/AK0Ie0JE
6SHqt9twTUC1vo8pGwv2dEtIEpWyW4hChQSW7ypsHaJKUOsZMsmjQOIFs8mUqNaU
XaepnvUn0wKwYz53rx8SMS75CYitRykwrsfGyyUA6GzkeuWj6Jt1FlW9gEBEqXbD
N7GDKYZaXZ6bWyCcUYWv0bUg9MkKI1ciOGhKiPTsxIHpFWhZs9eHh1nTzR+W5xki
6Djyr/J4olXgR7CiNboPMyDIzeBpqzBKVpFyBBCaMF+CKv9AzjQ5jBYw2xk+p6Vi
joOhmApC84wfujOZ1loP7jXiNB2kwqjq6sdUJ0dyWkWWjWn6e8ZDD1QHJtTr4qaA
Fg5IJIUYgbFTBpPIO+6e8NI59xVY3//UEEtY3wF1GHz9WVyi8frnpVl2Hfx4Z0PI
UF2jZi5zEfmH2XRPufC9ZeTebzd9f6sDqfX6WjYr3JHLd2xT2wRDZPg/u9+ZKQbH
8g2UCHyBc7lW6WsG2nwgahxm5auZ/0hQIT+GrhCAdecUfdmKtANBG21zcC8uCyaD
cBGKz8nFsM9iD644K05xiP/UcjPDWO9W5rcFcVQP9eZTV26VL9jkLgAVjwupPm2M
A0LWn8G0jzTF1nCKysG6Q/Yy10o83fNrVFqVuVAYVUoII62h+/V9k1Wr1H0DGaoi
j9k5xt3TbnMfVsHMbLQ4wU9CiSxwuIQVic6vfLZnWkXrAdaSvv03E3J71h817nJ+
zVeRFy2yAyBFW16qsYY8WMlL8Dm8aoIu+BHIXw9HDA82i4ePDuPFQ4DVYuXj9dJv
A2ZTgY39Vhf1ZqTXcg22M/bROqytb8xCQq60aPBWiJpDxssl8JaNeYsMlbT0jRZr
xijkj4w2OZbwVg6e83N+yXcVpsgsXY/PhHgLKMXwriwUg1+y7AE19Dc7tUSIonkY
bNaAJZ+aDa8wshFHeeDRL4IPKe0NDF/0PA+buc3TTV/brrGlII+swvLPvv3x9FI4
SjHpLp+TZMcB/gmo4V9AidKvULUuAmrPAqL6o1UHwFZg61cp5EGtuYt6BzUZgYtE
udsECC8ox8TsNwKALTHD63YyeFdMXMk65a9TtdreYn2mOLhiSwTAj/S+apMlDib9
CkDJIVUT3TEgrDiiglCk1GMZbbpYpTFHq98FF4DwJH7zOAC68/nf3RwrUPOHrPIU
Mo0hc8tA5N4uCfloi5pG0xrCgwwU5js1npaEGE0202SnCpq+xgSzm1SB1e4gj60w
zR1x2V2b/kwanLFs99tjeenCJMIASMiMtxjouxlvl1hUYu+/YwMXV2BuNoeiCsdX
URcJsHsBkAh8Nt3AuKq7WTnKpmSkr5DhEqugdIKJs7zAjHi/0XEgDBMlBxH/bMYV
6Ekefvvyv8h/dtwO0J7jdO37zLQTDY2UhrJPvs8/RS0+K5IYHmPqO0UVMMUCwt6t
AQ+7Du/YB+/NyhrQFkbPtmR+H4AVnoorSzKhsyZI55yLAfq1cMdXhqey/kFVD1Vn
OzjzrtwE5Q4Mkyaicp+AYLkQbUYbxaMPXWZQb1esVaOwc30/inSGulIT7D1rkA6s
PJEXAZnHwi3PttWhNzR14D8nEUdLOlFjBrP1VmdfzrNwDXYR4gw5vEW+Ut+9W5gJ
Dh0kgVMvBltQzaiwP80ixELl6FsP0sHezX+9daJpq9J5HMwIosCaqp+5iXGm3nkn
kqyWKIUBTB9bbsD/vgeZFUf1pBDs1JKplig9CiBWsW9cGxR5K75Ha9awC/o+c4Wc
0NFBhdC+xp67t6EgNnOHniygbkno47f13MNFzAaPpF9T2zqyjXD1sOdHCPsYbvep
lc0yWkaMJ3+kIoU3b3wd+kpBHm6L6mB8WXxemOAtorIqZCsFDUlc41VIGSUnhxBH
1g5VI5swgt+4nAO9kAl+l/SdpU4HvpEEkLLDV6wUbSJjZToyy6mYuuU+dK1/TjKs
qonZ1Kcxcd4hiYep0IgeURWkckEbSyvFGyWPsCyGYmOJhuN+DBM0QDPqW+v+qUVh
zwn4muWYPpiMd+a/CgzAUrA65J20ecsMt0YtGU3rSiX+3S7KstI1Q4QvnTXO6Fw0
fktY1pvIk2W6mmsSfiqCY9V0d93+W5w/V04pOmofzNELPj36ecwuIlRGgpCQP3IJ
9ewTiui6mB5UBrX2QLQmUmlGuJCPrf8Lf5fyaogmhVCj+7z4KGbn3zVCgfO8UwQe
nhr1TPzKFwfw7HKyPV9OOyTE6/5aT0OEZQbp5ySRU52L4W0Koc8TZs4W8EE13IEr
q7Ncl9XxMG7MEXRzL8QsBI5LsSknMVv8HztfKvctYnw/KbIPSTdBN3Dup0TOuLZV
DdWsPrHrnL5RRQ8sovuBLCS6pgCopVWSf8oKby5rD+mUO5VmDPP4PyNws8Io5nWR
wszhbCogJcl1FNTl+2pRxMWUZQcQ7hTy7yUlS03vvXiQ7/1LygVLYRfcn7lpTfxg
oHpkZzVjCRjyWJiX0IBrqwZdVWYZaLZTjPr2hjAlO08hEZCJEgk8IrAuRFcZKHBa
yC0QRNsGlxG+mKnA/JL9SEN9cIochbRhhpKiShiAPWWOKHl+pWiS+UiORaHdE6EU
J0yQJpmjbU2KP/pR4bmAh1TNFy8XULJBd9GnK0dIal/5YmznkYyHttWk/4X2s57z
oQtEXdRZRv721ZtUZz0EUivs6ZtGpuxMijVWXlQHD6dKC3ySqYVjysPIAeR44RhS
zcchdHzLdtk3+b6Aj0LRO27o3ZTH4nTKE+c3xfZon1jaEdDAlhIDGuNiGqRv22YP
sXWgpAo7fyboelpvUgSCw5sFlxedhwjpU6S4qV0bg4Hkd5wKxxgK4DcXDnedr2mE
eSENSFixDJxq25pN7kHLBO0oyRt/uR45rzWqKDj3wnlhei2nX9Bju5Qzf69gry19
IDyb7jrSnGkIVcRblcsjRMID5WqfFf1n7T2KTF6Ez6fHcmj99lEFhgEPes4d2S+x
+Lfa8bL6JmEt30E5sDLLSFslRvJ4SiNv2mCMhJ2ALQ05UbzC7npXnlj5n8aZVGnQ
zJvs/mVNStdKRhWUjnFLrbB6s//5BY6ruqYl7DIgeaCPZywoePtp4ZOOXDgKoptm
gIGc/Qe7YdPb+UZMGrMUw0D3HB+7KWWGzG8jFRowMObw5Ale+5RbR0nYp8llTc0m
8LLF4Tt0BBN0TahrvzbmyaiYFgvqABE/WlHTOxRmAdyN5jDiISqLQAlVPofynPVw
pb6bSXXHSMMe7PZzRFHlNBdKouJhGRsN2xAFdE1JLq+ugQrxmiANsEiA/J5h/aP1
WCxOFxFRs2Wcwxke60suvyb6kMWAVy7HxsGXs9ktQvkzDakBLOPc/Htq3sv/iAwL
EkU5LX8aNhTSZtpOH3brEGw4+6HrNniO8AND6cS0csmAYQfhYfnjiV8U0sYRS9wV
eDin8pLwmes3DmHYOuOhQKWufi8356GmjBLEAV6Sd8BH/9SdR1Qlmhd/hzVQgX1e
PLc7i6YTlhF2UJr0iHAqnMUdZx8g1VBaLPXrrHWJsGkSS9kIBZBuX7NNFF19j0w9
O7piFCxTXjC1K+21hLv9QSJQSoLjcOYFPQrUgSfdW+1C2JCad9aLHtuLf/jCCQoN
mW+MjQ1hoJ+v9FSxksCgPRWULOmap9nn/9ZVlJq6WvTUcgc0WtfBYcMQeZgmRi3e
o7oXvpCRIYeaD9H+nUkKWIeiczFQ2muaBBzZ2dNl8VsYSdSFzW0TxE38h8omcgsE
s/MHLjuRIfFf1bJg/s6jBn4EBAoYtp7JEY7W4ZIbc0ul5vXIHQ/KZbb+oOtDJS0U
2i38KIqqOli2hJ0kw6MqgHONEjrwtyi2OcfWlFSbZPzQhz2FLm4kw/tH8kCaX/oI
MR8BQb/jkJC2dWpkvfnmSe/EJF3OAusmP+EkWDe2RQ8IYhWr8d1GYPH0PsH3u/gl
bwamzdRvkqBcn54YD+RLsDRFIIUcayHvUO6csXB4lcOX/hR4dHx8k80SvNHyfWuR
KgeJTvPKVK6fs/Ogf4+iKS4kzVw4ymq1Os5Ch4w7VVjm/CCIXxgtysxkAcOcJdKb
ClcMinpzwxGHbE4nNp+SdcDaA7HzxQCva9jy2VC0qIkw0jOvVOGn7ODJv4zRQ8JR
n68TCOEhp9j+KRTeOD4ijTMuZgXcTsGmPm9vOBzHcCaa92gbBoFNHJOWtgsKWNC/
JlwztrZMk991zL8FhUgEpgVHMvPR3lQJb9AKin+C4WU5781joG/HkF4IjA54g3PK
C4fsCH+tUeqMhyrVZlymAeETIctA7f3SUSfKa1tXoCqd04UAVu7wU0jqWV9xMLI3
PAqG3LyE6o1Sp/L+0U977PSxd6nVENxwjtVoeagmBGKbbTroaneTGf3+xp5D3Hae
PbSQ5VZsDAyplS2s8Ct83f8ngfzmXJzrQnZWUFQ0zg0bNqTiKbqqlCbVtzRBc0zr
QNd7i0wni3a82ECg6bHxiVAULZ+iFGcQaXfXxnATarLxTtVWVfosOi738UXuc5Rj
Rrnktcu/q/bOgBSaU/m2DOm+yXeSV87xhxbupgZuwIMnaH7FhwPTrsw4GoDZ6Y6i
5YsL23U9OjmtHvdXwVIGVLEtmk87CvrQDI5XMd3RVs6zku5i5tx8XwZM/bzFYJAm
oM8DzTEtVD/F/4D86VE59megkgf02aKeQieTGHIDW+dcB6P3bCAgzMku1YOEy8Vj
quDB40nD4mgj0ymHtMIFiK4CDxvUr7Wo+RsxOAbfMcCiPPCr6FjQe95n2+06vxqF
MJwJwMRRMg8Y604LOd0X6Ir8Zs4r0JnU1NgTwUIBc/TvsCSQXW3hccZdMRbV9+of
O0lPJg6qJSA19o7RXD+AY+xzZKlMDKWDBgKox+Mt7cOFwtsHm5tMoKoPpAmN6CKO
Hd8QFNDMhwgZ2Iir4RV31FVqeSF0ywanTEXDOuTKTE2+lYNoN9KF6HC+YAV02nNa
RS7g9C5AMbwetuh4Qbir8DNI3UJQifemP68K8q7N/hSBtkSlZ1BvMvMuntCM07Oa
KhypTZlaxrJ6+crV9R8/B2Fb1J2xjchJZcjKy7t+iBkcFiNnDfeblaHtnaAjXLOl
vR/PnlAlj88oDGlrz6edHP/tYEpT7vglr2JaYJ0p4836lTEri8j6z1zKkVuI9l1Q
bJxNE1cGmM+Uc4cwz837uzyGSesgNgPauxb2SKmFvHWJA0cKAmR3cJ6f/d6dsf4L
y0pNoRc+UuRGNBsWrH0N+pyN0FmSg1VPoCTeiDaz3W+30cNjsDChPwIMScQtUaku
e60o8LZgIX8vaovRKJwjqPKvuNHhiIXxpRC7SSmGVcHKqEG7//JhCcHzarhuWbH2
0UlNwVRkpXnopopfeBUB/gSWrd9kOZlB/RpYRAqTTENu/zbBGaa5nQSOfJoBONmG
HTW5WRynNOUh5VRX4YUm9xVaeJpPD990N+++oN/k6QstxUc5VsFM0jd6JSSGIgem
dPr0aQ/bEFHRD+pxiof0l1uC3A8KFLKH13ju9VmDxo+c2BGYLPorjTgdt8zehA32
4Bq2BnOhNNKTjN3E9DIHe9jIWI0x+UBb2BDCuxCGpeadU+LIsw3fEaDWq7qGMoq8
dCviC8n5ljatEOx4f3VJpj3sI8hkMNieHDBe8xdR0dpzV107naxHeg6L6Qj0Yuvp
3sYaNCAQEeJXQcmGPT45bE5FS+Z2pu7OvF4mLcsrnJLoBJEqy6nLpN1vq71hkbyo
EZWYcYGLprprBSEVjTn5pU659jGZG5sx6JTmQRuml66SzZzoHN4fAT+viOxDDV0B
3ZSggoQd/9qAOnmjup+TQKLi1tUWIUWAP+HhDko160xiLlfmzLY30N67IZJpA+RQ
2riy/a853hCP414fmbiGRPQ1+rSVR47WHwL1xOFEkyf48y+hAIuqQQBUK4CquS9O
68K4rRXaLRVgAjyNmBKITxjvG2ztBDVLvOP8hlo8VwWvRx+cv6v3SQRm5wPtQEDr
SBVzNNG4kwZBIEbjtSwnkK4HGE47dyG5upNRlb+extprdYWp609fAmumcApUyJAR
jAHoX7lIyYSNWrn0HD6UY9/hZsZbaKp0bw6SaTTa0cSBV8BBY2Kn5BjFywZhCZ2Y
OXxSRdNSIVyYBCL3SeLmWZ3h5FNuKYKF52tzmGXBKP9SZ+sN9IVhasEK0UoU09gb
8ElHEA63rEBgR7BQ8CQDF0ULUc0seo5xn79BGCTsRpb/NmtoPu08AWJOJGvMLliG
LSsSzQ2lgVTBMJOZnKa9fo5Fx1VEyJGPzCGhCaPEY+shBlEIIl5KTiltYzUwRGNP
NcioQ0ZjV283FpetaWCsT/ve5ywp7IoKRoCF7m0vxlBIgJVTDcU+5dspGZWh3gXD
k5HFFuPR6rPpuY0AFbaJ3siwQMCOKVzaKCIPGRK1Nl166wUaf0KYFL5zWvt670n/
AdcKEBgHrJzkd0ZMQb3ACYOo66woYwW4AQfaEcWaB8Ksfn5nYY64neRUinLj+hOW
MDagyq00M4IkDRQiDeV0zns35ri7mKV4b0uko0Uvm1XoOCxkW/eK+AELJ8Oh6Xo5
aqCyxni4Et3+KIKXWmEVP5gVenlO7zhAx6VByL13wfRm6N3spUVAsHR7iy0ElCQ3
iiKt0L3xGGI6WHiBPHmxo/4UK8hGhJHJ8Oi0xh4DCmu4MnUuK18vlmR3SSn7skvZ
1bxsgYcpdYTvep0cUupMEK4UjRFYb/GgIoDwKKUzMDioAljhCd632mYAo6yYtwNw
JoksToZoqtiFONU2QDmDSZBLtA6OZHI0D0H9iYFBTJzRmn20tcClS9JI1sfqcQg5
FLMjbSp37PFRwKsNvluBlUWQH4cJDVJU5XpT12tw6HSBfrn+TfQ3mkwgZf/nXbGj
27W8W6YyrITqDN0SltbiNE8HvaC5VPQfyvnfsJGIJXELM1gzS6wso/k1wrhFLFvk
IG15fHsMaNE6hYE2UMDKzdQuC4eB0D4VBhd/R0bK3yjfHDwMCPU6dHefZ4cgTdn7
ATF4CFHBn2pI1aZ7LMq/yR+ZmWz0pqsm2kXbffNvku2A4FCkVLqGdBpQFK12kx/Q
ACKvfi+lFxBhf7GCmPKhjJAygZiCjHoz8EFdWNrrEKDlwvay3zj0Zca7e/ic6AYA
a1i3K7UTNOhl7Yrh2mVWcWbEwTjHd3l4Fa+flwwpBZfvNRAc/ipxXEPdAjIBEfjx
sTVCMZvCX/KPihBXikXydfzZcP1lno8q0kzrMDZHOPb009cgFRl7DyrMRaFpteAw
/VPqc8FqzoFmCmKrRO0+MYptHBoXSHbYy5Fzhyp/z8owm4DcFZjQDU4PLNziQ240
z3oiSXmJ++3pYzYgH8XfgxTgjzAvjPfi8IW8FxdYTAXa9BtvymXrSZzvIWmtpjAh
V9tv0VC822iR4552NlwlB/2BgiCgu4N+WpNx+iTbn7f0YxhbfAtSaapXZGzf9IH5
SDtjwG6S5l8DsIoX+88PTWt4dNERVU8nX2Q8JRwGXZZOdbcPsogGBtKccGcAbiza
a0VJpoOOci9JplTD2A+Dq3tDiDaIOe/bvdB8Z/LcTXWR5fUxiok2Qqt/q05zNi+d
aMnnIikmaBSGSEsPerOqYGcpGHeCXnQDtSUO6RsfzJhpC4ZX8UqofdvZYJcvuano
H+PkRV5s1onIgqwScer2L4Q4QjJwNesWhdm7n7XSqPtu76b7X9hd9ZXKX1ITokVe
QXIVY//jIhRd4d0rVN9CFvqv1fCrLJ3WiCM1FJFsFAJGBrimezOUURj2BC18yCZi
I+0xC8xwIE/nSvOYQKguW7r7BhfVjZPShltslsXxPlTHbm/eLjHK2QT4GECf9m0u
78bL195ual1zt2jrTZRDg0rh5SXoBUvvMktH+511gefIzXDBF9FIHhsY6+PYBNwy
s5zL0oCXrF6/wccmMdn5cOV/xWd3uTrRMVabpmuEy7lSqG3eYM1jE4Tjnd8/s9eh
/gwOCzc+Hys1FHzsbWvcZTJwRoycgX8xLknmRpZkXiiimUrdfiJODEuutj1D69C4
6BV52mjAC7eM1AzfKakKcsqvuP/LfEnl7pgL6VnOoK3/RK0bSOdDAp1gAzzp6XTs
h9bQ986sUD69I/ByfLs+1eVoIKC/+m3xAmun9sTmeLGLCIceA3sxxQMMAR2p+ypv
s0iqhgkHBDrlsvil5t0oPuIb9wCkIFfZq5ortIrFqbQbGIPgP4v0H7T7UNSgVJcl
lrOFYth0RNQlf3g4L1YeMxKY8NMHhN0JZtOevR83GCSwovOkQW9LG4iCEpSUMitR
KjdIPnMRVrpri+h4GLXVpQ2o7xht+5RnRTP1CdiNCNSykei4OXyX9ngt/QSdp99s
IjneZdHdyQJHvffvYZLQhaGjQJYR9QT9rH+vFyHX7Cy/KQjtkh1jPuGAmSRRWADt
xvrSHzAIjeAxlMTkMHrbtgm70NXdN2LyQXqMBJjsZa+GvhPJM1HzqRBOlofAc4rK
hzDwUoQ50aww1ocW9MJVuvBogGv73iked+mB4CH67qR+0aS83OgNHwfEmflvdpPX
tPkf9+G8VHxwmhNrrrrG/ZFDA6ODYMgHjuPsIGR+alR8rA46QQjVGP/BUaW1q1yJ
RR+7W1cvCi3eaeEgTUj6rUpfo7RV7GMxEIB2yu4zFHtIiDYIRGOnQS+/C7YLjhwC
cU3OOa/peAf8oa21arIpDqkA+A/89A0T7L9tTEy/Z8K7y7SdpGlDeuiH5LEYgMmm
013XUIqBV2oTHTnSbaU//ycvB2QZZwHSlrmVM6/Cq1EJ2173r9sHQmJqyfFAzjWh
YMzeSrXv5JbD0vdnf/YdTM0MiHvma1HfT+GpWBJ09Avnk0qZ3/LIjya5rGj3CPln
zyewk+tC1tSEd89GUtUPFcaEYE1D/GCeaKgqCwPAqo9dTlqm1xIZGZPsPYOuUG1A
Xg3M4uXdkRwJnOJgHtsGgIS50kNwXjFzrwH/Pn0N2mbNd2ZUgANV3muV8/KBjl8o
zOtIz2os1AG1BAv91Cm5kn4eJhPWlDybySs/LUkl8+r6MI/qETULWKG1DVKyKQrP
Z6IfkThBeDyN1rK3E/e7d2FJshBub1gwFErcyXzvxO6skn5WB+t3/YzOvHm0iN/5
eWoIHRBJPY9Q+tFKP3XgF9UoDsMJnYApBTcTce3wqYbV/CD+90PjIl1bpbAk+qkx
APkavKzC4MrOVk5vwAJTcfByUvLDmRSNv+XbhAbQ5P+guEQZ7UuZNB7ps9+byuWt
COC3uN0ubZKk2w27+996uhu0rS54iPpXej5cqZ3TDqp1AFhDTN5pqL4ZgeSSj1vE
OJMUDxeCJWdarxLRGWnbDx9gyrlw9ZE3uREdFm4K719Wv9SYzSy9OQ56C7pLYLL0
GyabyqPGKnAxzX04qtIVhJJEZwqoNagGiyRW5tdPXzdXnlU7TULhskuxce8y6Kby
oz66EZ0eQYgvduIkDq1ZPa+mL3qqodYjuM6rY60+h4RtQ6SrjQUpvZnNbCdrgaDH
bS+EVmNZ47sIoYCXu3bYddAauQJOfKoWu1yUT71F6qOPPMyxBcsrunuMPuQ+mW2d
sOE7Lmp8MWuznJCDJyp0BqjV2TlPz83qEUPjZ1xU67SuhqQkvraUOOl5dWNoSbb9
diRfz5tma4IF8urq6rpCoofiP5NdRstmBPu5A6Wc74XxRf18Ae+3J0hloFXKvyTR
CNXib++0FIoVS1L2bMkNKn6krIkgVhRxAUn7ZKW6EKhemtJLK4Lg3dOyKVlhep4z
2K2CSvRTQDAjJ+ObHY+foJOtDJEhNBVJWFDC0eSBt4TUI7X9h7arYUtJmtji0Ou3
E9iSQkqrwOrXPhRHXPQCt3FgttQGEf4mvyZzRdsARdllPCKcou2gUvHE9yu7hABd
vXZYwk8GG6JYCp24/XANxLmH9Sn/wMIhWnyOtkyr4TqC0y057JZ2YQeX85EPT7Ne
GD45NpMfJAFWLIYbcFewu4D928x+HixNPkX0iCEGgOWjuhyLjUfOrk5hlmhITPna
DJKrIsKen4qe4AtDmZ9vGX++VFGmgyRFl/Nj5GK+Ehiz8189gJn7VfsvcjAG8wmZ
/2zvlO7GHoImB/XcRGRJl7KSeKHceeiEdMnbbiLi6koTNM9RYtQVX6moxGx524Zu
dAHXhlSgO8cwWu3l5Zs9MtEKRjY/Mdo8I7YduH0jLGv7kaqUwxjljCQq2uNag3ux
U8Bv+qyAk9x2td+BzJeeXyFY84mG7rbPU0Qlra9LQuAqvS6k/EKqx+ZsSC+mwM5z
zYAcSVUt/lj/mdK+OksHPZFAe9XboVU1DEsV0a68pmBeV1bXnC1+q9gquCv+uAAi
SWpwvWYfkSx/Sbzzhvwnydg/OB3euMFhAYlPoaK0+6NmPmyWMLBinJPKscE3e5GR
ybR0Hf5fo1BQr0KwZqryaAlp3zJWxOqetvnZqvt2dOg3E1QXjSVY9N0btLcjR0MY
dulYt898YzQKDRTBUyQ7ptBkaO1N6ai3Ved4d6EeUowoFLroZ3pH4RCl9o8AMNq2
O4RdTJ2fb8t4Y6jBPHErDD/mbsZUk05vOsRSnPyEVUovWYNGcueAMy5aFsR6DWdc
4WTfJS+mB8XgB6Gswc/Zqfl7jN/RntPM4e5ry49YhVzaelTIDtJZm88iEZTjryTo
Qg20zH3LwQfvKVmWlvUnFqQRU13pnVNVx7ldJIog67papMaSrpH2uu7JVmfKbr8A
h3ivNZV7SxSHLYW6vweYqXrpcsaVvi1l198jkBhdpsGkK108aP3u7at4KBQqA6U+
p6y6aHHuQMhT7Uc0TSfRz0hU0JEyRCho5CkPo3ht7Y6ZHzLnvhruzVWILMaXe6Bk
BvQCtMFGLslS7Dkcfupmjhrvvae0I2YrcMxjHWul9nrwAjFM1s+dmRR5Gm7SHz1M
5dVgZQfgZdauIM44nAFx4Wx3BibNxfbhBQMAnC5WeF1vGM5//K4finqUzEj05WUD
618EsNyiHnXr/s77WwbOGeBcnow5HDWS0u07C+kxYHWR1KO8ArAshD3LLATgebVs
VeFpwZRE6Ntm3azEXhYnjUFlvrXiJ88h6hiy5SMhWrbYAazEnMdRR7KSJrEZwM23
pN1PEElmnjnp8WxXF7a9ldF3GW7P5zW3gDHDVQb8op3XtGHscF+87ujbf9fmKlkx
D0Q8Z+yQBIeK0GfSUSQ8S16zKEodvDfGTHY5CVOAjjm0G9JeKuttJ2SfC9EYNEYm
5J/jflKiQ2swbdkP2WomeIKUmO2xRL2Tf2xVNDjNmbJuockdMqr0hTnD/5wjYZbi
5qVXDo1NSz7qhsBnVVP+kINefEf4QE+7Xpqz/AGit520V/B4qJ7VzEIOBzYq53Jh
FBqvzTIfdiSqROogj1Uw7N80aYOjtvZajfNO4B5dOD8oZWR7Hn2mPZ9JKj5i0xiE
GRd8mkTqyoD0c2uqrdByhWHK5gMd+1q0J/21u6uf++F233/DGotxGxuZXjrLr+FP
1BmS5d0BuFTYz+RQBn+3EiI/6X05u09Db2huKHX5hNQkjrscBtWn8e67O0QYNOyQ
3fbM3xJFGPY/w1t8Lhg7h7DsOJr1BkSL4iGjOFmGYO/YD13HXN8qScyMS3Zb5Pv9
G8nK4iJuPeqQtCRJlNqV+74ECyBtn0IsJAjBJzmPskKNp5yeMYbtta6O1TDEIEAu
r6nfNoEd00dYlv0+OyGSiCcqJAHMrGa7s2sbloRISBGd4Q1SEKBdIsIfXLXRhtnw
bvcD26+e5q2jH19GOjHqKO+LWu1AIo27iPAt+kInV7TcoGpdNsj/dZk9a0T/FoDC
U/Tal1mMhBNlZX6S/7IynwZaXvD6a6kTE0wpciRoUc45nEdRHunVp0IRbqzyv3KO
pXtXdhFFd1EOwMSwKAqr94nmGUnYwCGTGZ4bowI/l8CDv/keynsQEt6G7tNjpibp
I7nBdO7vvd/g9G2+vH+P4mT6qmaihlJXGPleEwQzWfnzZguFWE+h1CXSoFfvbNKg
X/an7LP8zMan8XtoGhgdyfdGG0EpWJWyoumpASHusbgZl4KcK+ODm1+VFo2PGQR5
mISbvcH25h0fpZYiQLcdbr4RyawCs4QLtfwhzyAvY2U/3ww3YRqC6KHaMqRpxGz2
r89g2kk7RliIAUWJ9Ga+s3K0GexJu0wkVwfdFyGL/rY8Y1DUtP1dsMer9HL1j9xs
a7ZWU07Yf/slmrdJp7GCl3ibs7IcdPIL30g/iSRz6tVyUSZ8gkwFESc8j45GyTsU
Nw+C9SRsV4o59/ENjMs5MdcwaqPn5lfPCSv1rCpW0NWBf65c+QDQtnDRzHpkSebp
xKdqcBWSfyvc+1I1jgL2++P+8+8VDx2B8ETL5nCiz2U+SxMdXvMQ0DEaWTIDVN2U
3TxPIHm89I+tjsEos/bAMA7R3PMB51px/IgctX+eIaEcUFC8yW5cbEYhNEgbH/vY
7hqkUxwRZBGTZAPKEr/4KiOlzVuPW71k6NQ0QX167KQ+eUQAFEpE0T60UeE3WwOa
EYyQOJPs3zkh/nmsaisWLRryfJY39znALjLDd/yjoXbGrgMDCVlTKol7ZfS4WG7g
BQu9hVP60rzPEX65jvuo2Sz/8L1x4uyHLThA1QIc9DjbLlzROFrKZ7W6pcykJw54
Uy5MAzA0uJdiPXISaPT4HHqZkBYFR/vHkFtPJNeJaWaojnl6VQ1r2MXypxZDZGdx
RJwuaQ+LirR/f51cB78grt5XnV9SmCmP5oBw9vmNWK0I24xBhKI2CX+LJ8tqa8ix
ybNRYhyZcovzr0zQy659keqp1n7h8koFK0IlnZjEE+V4VnZaV1K4NuOdKbA+aGST
EYbgxdOewAA/TFFzw/h9emRlTBr1K2CTBgxadLx9+AlQsRO68umCtvXtA1/mnjgc
lGXnTeSvFOj1O9m8L6C7Kos7v5CZkAUmX/diRU2t1hOitUfLWiXO4a9u3V0QJga9
LajvXLsBvvi8L76TD/3EGsmGZ+jDrfT4eV/vpb1a2soos15w1yBoCeQxFTBVQFsW
P+EHL0aq7k3krYBDggTEtGFOETBmokRwAFTkVG2QgaQZNigj4gSlcQOp5H8fs9uL
MDYmGeQT6nEeSRM4Gi3X2+Nk5k0tfot0xmb4RhBqs7A07+20amroJsN1uxe5OVFN
gz99b61bAfJUkKMKVwA2IsbEzbU8JpmEpc0fKrFQ7LUgrYJX0bJVpLAmEKwhjCqQ
vzR9Ys5rpjBY9exG/vkF2RNaWyS+9JioL8vCUxC1ToWyve6d2dchc5rVMz6RzXaG
DgMM6D30lOLEMjeZQxOLYRoLaOzFK71OhFOkxrq+wKGwAd4ph0xdpmuh3TEeuq75
t+ZiC97mXqB75oY6haS2JZkrtqH+aVHi/yJ9KK1dp105WZnngqAeyDZDWpG8DBHX
rDsiK1ETZ/KI1h2GCh4iLdQmOFSTBhxEaa3uJi99QXdoUfK27GQQAHiduYrMdpnO
Y7Ic/BOcaYzNjB0khU0h/n6p7WH69uunSzUd/MX58S22Zaf/h8zBAEraKjkHoQMh
/NZsVlRSAVrXhA6Y8wTSCW7BdUflcN73HmljQ0TwFmdJh8eUqGUJ6fkfpEDnpTWm
Jhggyj6jWFbeve7gXc2SOPOf3HU5uKc1enN9DS3XVyO5YXocooDkd4C98nl0EeiS
gYGpbUjJEXYR4ALoF/q5tWVqP4wvv0vFcJ8lj0+DRhEB/GIkCJ2LtD99y3ymTt10
syK5iXLLHHWlINrOFM0dp3/s1HLXatQ1rGXSGdWjKn/kj2asEqtIW6Sz6WaySHWs
U9ngPrxHzy5SVhN23v1MfnDikkUuQkdX7VQRH0pWdp7AZKwzL1lr8mOD7IOQNboP
0spdDYwodr85iQRO5lNsVcIEZXGmBBJVPMxfl9N8kvtoMiN53iqGZIu3b3434iJI
LWKUTDgi2kn4eeuRgHm1UQKSpasnkOfrcEl9QMuWSBstcihiCcgkLg62JC3/PRdX
TvOUlvvqgpL3I1K5VIcX1AGLm0h+fb77H56H5tdlzAdRCe/5jMFcK90oYEU2cz/r
qnjf/ixGVThs2AJC7Oy/ijrtrePmJV2NO5OZVqJRbKR7JCwlzrE48FDafR+oiFaY
r4reuEThMfOId6xQiMkkM23LYBM1zuAWwKtl0X8cbGqF8wEbbISRtyJWo6/7Ul9C
vy1UGe109Odxtd7yHp9PStFT0A65I6azyeIk0jVX8NwRWcFSZ+wISMMn2V7f2Ss6
qEigIdR4S2kivJKRW5GGEOxlZsuPQ1wnUxxV6rgM1Ww9UUfIoUEG1MItN0DLg3y4
aoUIY1v0MZOleN9YNJZVpDQkLkSKp33OyLsKfTEZB83XzkOanqC2on4fDeWXE5mK
52CM/XULN9D+Ie6w+l2Wvqk/wLaAqme5UhfuaSIm8pHgzW4mgl42BGXzOahd9sVe
3JQMTlDLKBzf5SDebhxDrAOMK0XYABATw5w3LzvDQLpTqnbL3yJNxtfqcVYoi/NG
52yPeWqd/Knjcjqe09rHXvEltspEvDami5AkXYMW1Hd8GquzeH4p64jjK/ttHvKS
t4AbfqyLpBcSUVRtU8LdmOejd6QF3I7F3U6NdPpZtrFei52de4pCgn2cq3Hv3q7J
2ewQTXp5CafADRNWj9fPpWpddR0WQnfe7U9LXxvFcuXnTxr8Gof/7tq54FQd8iK+
J9dlsXwZzeR842htiU8rwgbl7l8mzDH208cOejcrGt1wKIwjuIvnE1UTgu7HmNvf
hxwF81KsTgSNJK76hrFZIUZNAtDIch0reuAcFFoSV2PxF+u64/KeI1dwTaZZ9n7p
zqa4f4Ok335/EPdahRB7VUSmEiem+BwMxKHpqApeNmxD9tYxZLuw8A1vQVJSNdz+
LJQ+uV+xvY99vtBma4lHa4GgBbZu4s0lMvxqMJ7dfFL54cu/3ECw9itT/fSo13G2
DavS9I34rSuILjIecIGPK4iuT6iMQR0/hVjwkQZ6giqtfHX71/ikZVxBDVlyrMG/
d+Z0Lbqf7qV4cHelrpgKhJ3fxbhrGNdMqAVOHQHdnIS44sKkoGcm2K0ds5qQ2rcx
o5fnPUdocJShnmPYX+8zkKQjYpxkkKsmZSlblesKJ3baZYk2fO1Lk9C68zxkJch8
5cPikANZpvnx09dSC2z7Nm6rDKfs8s+1Hlj4jjGrlf1Sgpo87vN3kNI8fZfnbVoh
AKpvAtpgWwemYhTQckn+BdIrvRrtg+x0drpwl1J1cCzbcNJ5F4k18pIsT324Xl/0
2YmnNeAM5rMXagpSGdF3+34o+vUlvcUOqN0AH2DHUJjeDYzLc0PqggRkUNB6sZ6x
zpR52HFy0J+Cqht2syZM1CsKV3dkTe6fKW0HHToNzIrHka9ROH3yT9iHpzz3GMLJ
1/4WIZDI45SId4WEesEdIDAUPORpe//NhCcJ5Ch3MfFgpBgbj+1wdr37IQf0EoMT
E39rOXpayj4jEjcd/rPJlD+da2a07RwqnWkmbQWYSiiSgBS4Cm+gyIEaQbf1gKYp
tAs915+OfgHey9Y5Vxe+U0HJEeweSr6MO99xK+FHP1zOtkfhQbHZttA21vtO316F
CsDZ5jGhs+CkjxooOKmfMYBadZ3VFhaLKJQodhGLkrfHmeUyLtNyskBeoecWGYjG
v8FSyKLpg6jgoYP7Qd7V3TRAytxAPyUy91G1rG0FimiPvmv95gLX8E7yUnPnFBeE
SnRGS/ZpVON2YrDyFWEKepBKZc9SaNI5s/OLpHQPffGBbJ9PWXOlOoDQlzLJ8Vaa
x7Klf+drioBhBxhnF11qG3+ZYQBXSkDAaJj/MSsN7D+e42QszA4rgU+v25xGRgS4
Jhp9tyPYnlYD5FfYAHWMNtORtPnfH/Z3Vo/bGCpQoefxLe2CywB41vG5IxFhIrMq
aI8G7gZwSRzVhmMQvlKjMc8E9iMyVvXReUusBgraGsAHg1gD5p7ZSgNh/gPN6AkP
JD2KYIM4l3TyDfM0YJTKO0a242QgH56+UB0JC3Q+j+vegX1Qi7Lr1dWoetjtmJMy
zsnyZuMnLq7PeoMk1FNJml32QCmHUrvZc8imqr4mHXbNh+2crNkODe2UemJJmdg/
nzRifD9XqWYrbrVlDa8oal03BRvkQvTZ0ccJ/eDtkYuRAiYBIYy15XvA+KijwTCN
s8TsPv9WN/Bm5lRV2sx7IHE2nkDsDbvxo/O5m+6Ibp8cz5ldrU8eiigi871hJy7R
niN4xVkl3b/5QP9+Tf/JRnI3y+ILS47UdfAQxm8Ym9ixs3i4eF71e9EjK+kFYzW1
j7QqPNJOXjCoO4oQlivabPqi2JqLArMzkRphNrxBsb3diwU9d4KR+9xInDBS7WLi
L+D4t1S4q6B3Gl2lP/+Z0oXQw11DuulM3sK5PoF25xTL0XXcsj+xZXVTn2By3M7y
NbYz+kfF5/tdXTsbKd1YgzOaf2RCYYEMxdD8m+ktcshVsY55GxqjFHeSTzf7ruM9
REKQ+75WI7TKvqGNRPGrdsi5GmHVAQjAt7aTj0rWkAdgVYXpEMgizeW1/NTeurUJ
9+WBaLfaKwYfC53HQ6BwfAcKGx4IXU7z1hT6L120LHGctEKdRbc73Qq4h1bH+olA
Gd7+13KyIw9mg/xD54LUTtNa6K9bKjP+uj/pv0vr2RMXLtXzFVsUMcUizHt0OP7b
NJ/OeQLWXXCUfo9tp/Higz48JoANm96gY4Jfztp5p0lIXMQ6doN1JXn3shGfA22G
7PTxhTjkN9+lZi75Q9ZWaErzMhm+nFjDNFLVwKmLo6/SfLhHCXqslZ0i3Ws6t63i
81HbGGU+EQmW4lIBL0Ld68J2K3lwGp7P7iqOWpcdOYgLqlEoNeAPqveOlBgg5reg
V4U7nuKczFrXmofcfiHc7YqhcheSF/tiqIeM3a0iKB226DUyCjfjhYhnsf8skdfK
cKt6is2T0VLgdblt59EwKyyaqFZ9COif4ib/TmXPHdtTfwbA4Rzs/naofOhHWWml
Knqj5HUkr9Gnkn0u9kQzBybcd72r8tMDlkGmwSvI2+DyxTuetL6AMX5LaS8nCzzB
gSaly8mUqvlpXk9lTlWaKKlRFoNAp9NO0GryV190CHSAXHNDQZp9AGoTPnp7RxDX
U7I3wF2xSqTR7jbhgK9aZXpxM1XTc9KnBb0rEygRJFXp1OAT2azXFmALwLyqRHiS
H69sckk/SRzVYUyMXUS1ZM+Z6siLAQhY4C38bu+gGfnUehOkFkjzUIEdfUN3Dm8Q
dMVJLDbsA1DLRRl+0b6k9p4+h3HJSvaVY88xlqtY7QgN2VquSLu/zFt7GKh7VkAy
tjItblTZZ4KDDYV1SahEFfd0YU0QcfnQmDTOB5s4n3FERrXVtGR4w1eR/+JXoE2s
Ljdtn0ha54OH5i5tpTccpUKnctQLM34rS7ozpmk7S+hiTcLgqKGnTnP0FsEXVdLp
JxSHwiE8eLammsPffEyWgEX4vErZmGw6PrG7aJyB12NF+Ss/RDfGsflkwqxxOCQE
Q68rjS0g7r2mHTo+cXfNl6ZzXvW8cT4TXIbXSvZlLBP8HcbnAbSUYGq+2QeRn7iv
NapY4IVcxt70Sy5kRXqfs2cuvE3SMv79i4/1cDWz8INVa002nuubvy34TOl0MkPF
xaxXVms0/yzNASGSOai1bCRyQanuaJkc5oH2jKKVpONjvtE/6u29p7mnnNukGlc7
MAbFIRyCm2Ywhg7//llQ383TGKA+AYJFostTFzSM+hfywCg7kDQ/zZ0aXhprGnYv
+CVtr4bgNJeOzlpcGwf+ikFiDTL2RGh/Lpm0s+KECUBL/6kMc8nlrYLXKav/0+Fs
ccQgnBodA6ScrAl8qiO/Jt2OdnMt7/Bv8DheXumnanS8cOf8hr9L5JrcztmIrsAg
mqyEZBjMVFUttB/b44JaLr9e/l2Vw3t5LbGL5j6OSh0JNbqnp6YeFz7e3AyS+oaY
4Mymv5o8zNBewq+ccXVf4NjyvT0LyeeU6RH9C9AaIT2ioFb+Wav9I+7s9ABl16gl
IKGoFOy8bDRNAd6lpo3fezABCg/I2CGF3lqfkjPi0kTP3r6ZC51eq4NV1xg+Chy2
4EmIP05tdKpdEonsaGRI2hsONkv5o2DdVtR+qpSHNfwAguNjMEzv4aiDLjQvX35x
iYcFI0Dro/v5t9ytOuWdLBbbS/G1tBa7xhpnseo61YMiU/eYH1qkRy0us+6dofh0
HvqItvPoyh8YbsztWcuZbuCvQ0vz5p/xGNB6i6Y3LcIfxvqfJ75qsOZnyoKrv0gc
hEvw+kk/JgiwJfBSgtRFVi2xOF+Trpxk+E3uSGVwI9MwiDepqmi3EAM6NN/h+ajK
ZfpC+yw9oq+tWQ//BZ+s/YjSuwzYKMI1XjwjSahtMyHvjppenVceyn5sYtjb7b32
658zwwkUm7nT8G86VHnCv96pw9kEa4JnbkcrXv0ODmtvs2BudtZie/S0szNDz3Pg
mNdXt1tQhIovRGU2TQNdFSD4qH8ZKM2Bph307FK+VimaTb9KnYbd0I8DfEHuzr+/
CITCPtCLQfpNvcKfToVQNs+FVaw/FMNKEWidfZSkns3YKBIbEecvAqsyoTDHx5xY
0VvfFCG42Nr61lD0qkQfhKR6VJPYhth9VjY37j4qGDzOfLFd0IPCKgVhviRyC8TB
Z4EDMgqktbZXutqZOTItWbf9hefCtPI7w0VVp3EBm6Qr+Y0jHHzG8se0E3AHHCCl
6lDLU27k/5VAV0hbGlydxVMzvvTj2jTy89uaygpBh8O54TmDN/rX8iOySSNjTy9T
dNyLp4D8WRd8cXL/UIC4wpq0NvIAZpTjqGeEUhIaindQtYMafeTh5WNLOx0ZxyTY
G3z6Ld2krsWMMS+4jJkURRo26lYnvxpQHL84A5Umd/LhB6Rp3UMt5kTDH7uHUMIk
ON5kptUKSDYaoIu0fnI6nmso6Ddis/C3wu6ANrr7qcQ98wgY4whViv2md5av5WDP
DCBpkvYqj61DN6nMNldHRtTSZhW0XR2xuvIswz6KWmVQE+8WAmqfY9FlSSVaU0j8
kJPtwefAkdGepgOBP3qocvsbxweAYrpT2se00SKC1bxUQkrG2EZiTcdzM0NiKFEP
gEMiw9t+ItX948BpPmR4PhAHXAbpmRx8BuTUG1Dn/UL5lPBfDhW82odCrm8Mr96l
lMYjD4Wo7AygS4CY+0r8oaQzd+DjEb9/IIJLEo/NDMggpIiIEO9ktos7ELOOGkK4
nH0dCg59TIJ/DYOQR68A5S8nqesJaIOoLubLi2w2joRgfJs+vSCNGOtCNjZjQdIU
7abBrB6AHNkuF3iuRCO9dgq92llIGB5qb7nX3Q5tojdJweCoKN/FfndEjRkCpxfY
1VMqeZAZZOs6IQbJXDVS/NcPQnd9rP4StYpgyj4EnSpJ1h/ksF3SB4L0TRJdixIy
tdmvsyKGw614tBpGHKzNCNRZ4nW4qMlVFKMHeEIXzq5AlZAp1gjy4XLJ7Fi+fJpj
wK1gu5efGr7EZ1xF3Q5qMMDpWynfKztihU7AyV/2PWWnZcPbfLDu+dB1pZ+fdRoq
pB4xR13arfnSzrmx9yvBRG4AUBfpmNRGv2SyQAiIZuo7wB2pChuD4O5ooes0yWpN
X9KwmtNO2CU8pEq7MjC3RXl8SE+eketewOeoIH7cRVtTdkVDaPEI+1CTwC5WKqM/
N8mW5fd1usTygTBZJ+fY2RBo6RvSA7+IEw0zA9TAIF9nPWvf75ZHxnf2NcjksHYR
ch45FtGWzSc9Mm1ukc/GD6+RoHhWR9g0NixoFAce5HIlwdDaQEWfdjhVuRHpGEwQ
/JSubnOb8tjOcf5BxFNBXaIXhxE0B7fxxducAPvM+IzMufIhier6UXWjoVUlYXha
+FYHTrwGs2QXwxmS/ncV2qmnejvyuONwmMd/BSQLvRJeMbM7IXSO4yvoI4EnPE5t
pfaT6APIEzbzAzzspoOxaOedq+2u7oGQ8uVecHU8no4SyPeLNaylMGNm6laZta8X
htk2HBaWM2jmYQ7WGtau6uTTyoUH9czuTZis7vfBZTxxlyv0i6AnYaCk5+muRcRx
pSHdQKG8E2C4Iq9YBlQZLlul2lNn4aEm2GHyaEOSLypFgwuBgp2a8sM/Ao4+867j
Ba0Hvq0zu4rsLZRkP4gJEX92c2KzPvgLAXLo3xQ8eHt5cIJE8n5jLUm1BCKo8CMz
8bTbxmhpVuZ3SJEbTgIAP/RzIlaXfMOzH1W8l5Fm9cEDD5AdIhxCYbYC7iM1ftq4
a38fVl+db1wX/mRCGrffY68vCkZ0+LbrQe/bl/EasHOSlejA7kbz4y0f0aeqZiCb
rRA0RuXH/Lp9UUjlvzOzKsZ4iPj21FYj4BHP7H0hE/3EjcFHx43A5aC2GVOStR9t
FobE4jFJvluEw6V8+gmVmH0nqmpua+UbgvuNEPdwO/aAuLKzQHegeh9noNZYu0yk
vpzdeEvsYh1jvcwm9HhnD0kfz1Y462JpdWIjfjC36wkZhhncx2PKwJOBuhyTDPCm
n2MWVQA7d5wc57rRjiCu870mm6SwmgDIe1ze+2kpY53YKPNwvTB41IlB3OcsD1kJ
QWDA6yPUCVsN9/Wf/j0YmnRY7olVce0CR1RIU2ZOV6PI+ZVqw+ZvlXIwcjdHvth/
VeubbLylhTEe2m+Fz8FFdGaeu4kcSAoTp0njauiqeHad9ZBOiPyUOPAsOTIOEQMY
eYoHWKpJwhJhq7zF3fVOgdu5HF5iRD1j4LUD6C137Zun7WkXF0OwLACjNreB/lzt
VUG3EEAtSwQzu7IMFtKm2gvp0NQOOlPiuTKOJiSjZqBFoIUUWbB0hKEuAHrmKGeP
nvYpRQHqQ0HvZe7PNGC2CXIizDeIwyKy3y9Qd0+ys0Iw55X6tvsPGnoRFSMwy0FM
EW3OM/S+ZWiVAQ+7u0j9a87+DBvxtAtGQeglQiZuxjYU6q3DBcJX2S4wNJW/gzAx
hG4Rh4JatTY+Mwc5YvRSbXwWboPIMUNoe0Vb4kSN6cmKZhnRyH0eM1umx/BJWVH3
xZthdb5eGRvJ8FTm1ms2/za5OeFfGDgVbkk1+nSsQuM/mjVKGJdPu/hRc8VpjPXf
3GbYFxn2MYkOwnXjwsrBNRt56M29sycJm/hPWVS8X0FZSgT4CpPeGm/kdMHhzGRx
ruu9e+VS0iqanJz6zXRIAAzlRzrWqLQE54GKZxOvNwSjuWB3nKyAwNN5bvTvKZq+
4LiM5uS/0I5pPWWvTxElANHjwzazGKqgGYjwqVuCuI0eHuuUZJ3fhzr7CfLvnHxC
BWcGfOW3Pj7vvnuxHAoKXi84WRtw1tXoyp4MNneNLTmzdwj69mxawYRcWo9oiq/q
x7l+XKFCApnwxXdIU1McF2vQfXvOXHl0QvvLR0ZKGVkVongOi9e6DCv/d0Vjz6B+
U6SsD4Q8PDbKDYKBrd1Lg2rywE2wwtQGVULA542UipDRnry7D+biGJhH6uKDyVGJ
LidY/bwz13iutS0Fw7NFw1b3ESZb3mjjG+W53sANsOljIMTY0PvEgND+PJQsxMjm
iM8N7TCmOUfys9criSXxEDjm1Uj5KNC1U5vH9JHjjL8NggD9qeRyBtKBhBDv3cwQ
HYJoDJtn6s4nq6fLDB/5QKI4UlKtep4+iOvAcgbf+peVyJwCJEEwK0hSXp8Ea2DF
t1yOZousOttSqEIy2VzRduv0lTH10utKan+YfAUMFvNGOoBK9yq6/Roibbp3C5od
BQjvG0ezU/xAbQltOxXLzImUxcLqSU/1DPL2bTQCOq1JSM6x0qGjtfGp99gm+lxB
bpdpDEpOWkcq6Wr/Kk2qUcdMoDYSwRNwYhMzDy4yn8NgpXl7Zd7h64ZKMd/spfxq
wjyZlWGP0q7r3FdbXYoPhAf+7FFIpxj5S2ayQU/2YeWvhnsR4n492dS3hwj2KvfZ
Y4Vlz8zwwIRTDejO9gDIjnK5XWNvyex3/9gG9Fxx+gsYinLN3Zzw1uOUatBh5YqB
mpG3aEKLUooBKHiUO3Gf4L9Nd3+YM6JojcDujp/0gWywqYE2fQc1M9mkZWa2Oq76
2Lx6+rzCIc7IEXpEto7t47up0Nl70V+JYPpPp1oZl9pW+OKaZQrYvp+cOotPK+JI
oVI9gKW2XEacWDxpd1VB6EnrMOrWWPhWOine56+7vhobwApRDy1A/qJlYaAAktUD
6lgAOWxs0OEATwcPDNshhDKfnmHFciJIyW2B0Tt+MngbVBpZzgNHMY6XsR2b6k3P
vOMW1y95Lpoq71SdIFyDa+aqhMil/SMrArFTgZGRSjGIuamCKyzSlbfTwVrTQGnC
4ZPwYlbN88SSDfh5lQUe6v8VT6zdBMjmDllQCFehJhP988V77fvPtinC+NDhWG/a
E3Zj1iaa6p8qRqqJk4PWEcuMG51zC9YuHbRR1x0cVdTW8Ob4MGyxZ8HdY36jIWZn
NyOAGzLTgeGUEx3/Y9323ljuFZCFjuRrWhSOj3xApOVmOqbcV/n7RWzVaLwnD4D/
sb0pRfskyZmavilekBOHVCGlDnJoYyO0M/lJQqmSmyvd8jVwMA6BmpaVJaR0w4uT
XgHnVgbZDiv7kOqUoihchCXQpZx0+kL4rTQv43TgJDVOVe5NoGFqiLw+zC+OeGIV
yxHhn8NXx90/v3gRAyZze62xemiAzYV+f+vahhsu6agTe4NTwd1R++Y9rF0nPQU2
aHJqpj3vpqbr+fZd1iWQ1PzUYQVjnY+GOqemlM1ygt2Mvr8xpTLFWSBoEYfAD9qM
uB9jwhJfzpTNer0tUdsXKL3dJNqooyaRF5rcrKEMV94fpJR8fqzRhUDkS0wlQmsn
TK5sRAPW6G55WpIk2QdCEswcx7XpTgO8EfLNfExBfnMRXsuSDqFEEXhNz9sUyJWT
5RmjgcmTRd3wIlcASIGlMImVbNthS540zxRHnkFZQD61wClktF46GuGVUEq3N/0t
tw2dpkfdSgRlJSwtr/h0dmasKKV0s241lkrfZE9rVfV5N4zB+wGgwzgqyk8XQO49
Px6s4XN9lZmoQted9JdqaK3qu0RXsl/hoSzhRQRSYe/fmmMz1eeRh7rmr9AC9CeV
W0wP7ZzmoJcIKYREDW34sB/XW3Yvfr2vrQ8r8He5m7pL+ZG1WwoyFUc5yWdfLgxG
C47h123TWXdfh7hhVS2Q3SBrkGg7w90mn02EcUMe4fRiCP6YcVDj5Os/vqEqJ06p
6sgtknRZ+5MM/2N2taflghQqk1vR6hz6STdIJfOwWa/EY6cG7pYwZ8yLHwHNeTLz
CtRZ76tuNmHewQeDeppYeSnKzy2TLFZW4KpjrSFt2Ey2ujkjLByLAqs6SSlS+fHU
1vQeYPKALaefghUzE6x0Nr0ZnzD+Oj2xpEWEZzkFFvx2ONnrFz0+tMIzfQ6Iab0y
VG0jhsJdNmTGInT17Os64s+dnpv9hh0UKnGgMuBZJUTwxTF9QE4/fV3t9cC9kXGn
i3mhqZ8rwKEGNJe7SmBA0CYrnMSeIeSdh9+a4E8duiwSbgs/W2fk7a7Om3Ne6wsB
406NaIJuYfae1eH/qnv4z/Fm6d1LV+t0GKfM/siM88fSgcMIrqN4p1C1aeG+pvAs
Hfx4qNUzU5vDyXMGLVWbnC3qzmKczKvxB4G77XHqw2YRRzYSJH/OVRLIZ53L4cLh
Cd6AHaF7722/DvhO+mmB62pC3iBbaWgX6rhkN0/hsz5jjeLjmGs6XDfqkebI/n+w
qheP4bSSpf5H34O/qfREu1d0aTmz7+GBVlwQgzQ7kGvbgypHioY/OpKc3YqC/eOJ
IS0Q0gyHQf68aO4LIp4prGIMSN3DVVehim+ZT7Z4lY5y67AxoAfZxbPy1wcRgxLe
xPDFGPyKm/R966rpO+tkgLBpQZX6MxzX8aGOV6xQuz1l8fX92XCiG1pjSrFQT6bX
j3K26Osql5kmdTLZBCw6L1lzNBWVpe/h6npg50OIt8jijPwXFVdRdYERlCooBCyy
J4OASeFTYABVlxYBBQu4Z+iumlpMjl2nYtZEsAjpt2E9dkxnZYMq4DQp3US2xPza
W6Lphf5wv+V+A5udlLkxMreGxF7KKxXDhFKDQVKb5U3b4OgCqx6e7CnU4/4PJX+A
5ChZsVe9eoFK9X77FlUYl1Nuao4ByFhI4rtwIBEVU+A5i4R7nxJCCfsw/d6CUvtD
V61BEVywbFMLrSULpbUtM6tFwr+BaOy4lWNnU5x/al0ZxYq+JXHWDGTmZ5JpzyQD
AMzY7pIn2n5xb+Hl9X4NWGYBywMXXbXcmvaoCfFGxc1/kwB+FsW+AZm3T0hA8zIs
ADfW0Q05hvTYSoBvc/HjuOCy3dRDpXT17YtUX72S8WKYtq6M80ZehkSRLH3+IJ2l
DuSEAi6oYleuopihGSPVmSDmnNMh98TEtNwn0ucfcqa5TqEiolqx/owVuoY6X7hD
xac/ORyNP/oFV5/aqWZmyZwH0F/Wg3HgOpFsaJa9YImWzoblTBg6yqIkKAa7VIPw
WwrJv3vd7NR3wky4Ag8+jYa95qkOFF8fg1Hb/EIQ9FEP7Ox/oMg0ZPv7FoZOgCkP
srtwkGaFm2m/iI8bPSuGHoMyMqVQYjAQwBMvGguzoUF5c8lL2W4Xu9q63sMySpU4
pkMpz0LzNqZ4XEIuR6SrP/1IxkauQZkREyF69HfknHZiIFiYq3+bL+sb8OykJtmD
fSrRArkIlr0JSMcXEXvT5vtLuphUSj5mB0llkoyFm1mA2fyn+3oQ1UjUaGiSj2I9
FzebIJjLuyAqGtVqwL88NBC3cGx/PwekuE0uik/09YH++9Jdywrga/S7KQHCwgf5
ROALDjxbDpCxxbSVCFxiVnq6NWW3BUhzPOZGI9rcVvQkw5hyiYVHLIC4IUNjhzzo
A4lZ1lPjJamqSI0/FVg3+9gCyciDf71HCwdGQXWThANt29kVozbltvoJB3CtMMVN
wXRGjdwQplyXof6hdRXzUpYrY+u8idueAu7/91Jy37dWYBnmQGEoMj2ehRspfYjI
gY+hIKRGA0VymGM9y1D81t6YosUOX0RUJabr0j3Crati3g7mXPPWzJTgjpk3o+OI
Hpx5xJsjzcqVZOKRwtya3aYlPtISbxZE32Fh+ShRsY63mLAbBcyd+q0A6u4MqqKM
FUUx/JLj/UGBiijeCkRzMNaX0shjikFbd0QWg8FB8Ut8z+uUo4sjUbgWosLPq+Nv
l8Wi4NHMMoO6HEFBSFFYfvX1Ci+JflmUjWj4AMgJxJPqm6DngC8dAVx+r4Gd4ey9
V5ec2J/isdIZoYn6UhNFwFrX4+Yo0Tu97Q6i2vWu9nOEOtl2bBLV9kd6bb46RWJX
BnLk5TLrjhNpAyyqOw3q0cD4JOSFyNy+1pzBUpY24VtsEtWnWV90oUtogpU6HAJj
KVnnj7WHq8XdFP/44hmmXQkeNe0fJXQhU7PG2jvNT4kdftTPjg7ACkvMLKJf77Fz
U6/K1rEuUAFhA+KekmZX7EEfC0504jE0+kYaBk2Ixr4BzSMCvrXQ9TqPwgzmcSPK
ssS1v4UvXRIpjeRmvicWuu77ijeqC24HRKoZ826IJcQU1sW6ehtt7/K16/fuzMvn
br3ZbLkuCJrAUx+6iwkSP2+xDIkjrTTcG43i2XpTO3zffhLKqv1GBfNBouLdB8zY
lKKtiMqPVw9I9UIEdD0L8XtDUDBZx0PFUj43O1n9SAmuDUIB8xVdJ2KkN6LjoI1r
VjC1XXaoziL44WtWvzzUKxjMCJh6n5I5JTr143K+YVdLN0kvLmLZcAIe35Xr4C8N
B1e/qIkcuUqe/RCHofCAHz/SWjwnjQm+1MjwCSjtyxj0dZVJL1B0sRJIN9McCP/H
73jG/XirnVrGOU3vXYctg45JdRgDR+NLRV4mUlzfM/jdR/JSGAS8XC8Iexw7om+4
6Vv/23yUaztYEm7rXZVsVvJG4CA5pPLtAhHfh2XJft1QPdQ9JNMoZ3V4XNk7nmne
ZL92retJN/MSj5Jgpl5ANYsodNK44Nk7oCBii1ZWz42TvdICrDBEO5Fps1aeIQj3
qHlhnGiYd8bQ0wEOllyq3kNAFPcaaF2I+KWkC5Av9uWl5Q1uxGRiu9xNqch2Nz4A
13GEldG7WQjM2d7AVQxArQjPFsJSSDs7djRXzqXM6F4vYOj7mWiNvzfmaaTPUITk
/owOt2uDR6Uy3UIlzjt3dCTyLKJr5WdDWYAcMYF/krBCJhNbrHQlbrMDTr6V8F7o
ugyjvdnzbJ8+GaTCXXAATg5J/ixaip5IDv89SJz2BEwFBit2aLfUUtaqE3xid3dM
vAzAGl/XC1g3+F7/Y0nSZeHOTZPnTDhBjKyAioCwxgEhXLBMf49hfEgaUs3PFH0j
qlk6ELovuT2+0S8yzTj1Nry50J6jugjl6T4ZPqH21lBiy7md5JYWVfPSE7BrGdLu
evllA0htwzzLLWqPmVgIxCEGD9SsJEOi9RKzCXpZ+z0F1q7lI2365Fs1GhqN54j1
lK6M5zHhFHEAjqZiwXwhJHXjUiILldSifK8H7rs/n/yuaO+5EEtb/eBo8MK5xkLH
6jxU5nhnGhgmbUX44cBvnqhr5sq+LkMm7zuD9zSJ6ZMh5AWkQAWjQztX2Kf9sraI
ZJfv3ADN+DDl+lsw6tLwrsEwDUTBNHyjbk8YvE9xAzqLIr9MciFWfO1TkCylT4Ec
csLdyojcC3tJI9x+ESctPFvMaIjHj1FO8Q4xhng4okdLSrsTitH+c/Bm+tDyigiy
qdHQNbP5iFUy1FlLx9JT3O+60SRJWkxOQxrgVs8yPOglhwfh/369ECGrD7KQt+YB
lb38+K3PJDRX3l8Q2OmIVoeFZDak8CwTV9gnMF/thML/lmAh2Os+4VKv0UnP15hm
m7PfzbGa+eB8qKJtnZbUtQJxbsss0NnGRJHNHRUxh0VxJlDMW8bZyH6v1yU2r8cQ
JEvSf/BT/zRaOuIAmPmGo2EO/Lm7YBxYGBTUga3qizXGgnHL6LD+QQPbBcQbW80Z
pMZdlLfxRmE9o5IG43gu9wDZtxYdtcRH11W0CtZy60FYcQTK1Gk9TGoaaKbly/p8
Kj4uuKZzCj/j8RSVSpohJQKsaULSSHNUJGhPE57R4MwxJfof1Ps9jfPaMWN0rJtF
hHQkvnUio2DeZvuBsJ4YkFp3mU0doEhNt7lxpEnuSBSmhYob69VDHakoxTJFg75k
r6GscStEAarcxRHqUqycE1kn2k97JnmxvZ8qiu6dIjM64jT9RPsPmqBwj1Yv8ZXE
sQd6gtJDcWcPnsBf7Pipxl3TRYQfIQN3otBQ4u9Y1HzZJBPdzRenUAi/ms9UbFQp
HbinGopC1Aiv6LgRj9SDQzD7MGcAm8ihGs7SjV6tFfvRG9ubp+2onJJYh5K73Rw5
ROKUvLyNCUm8CI2eWvAAJAy+139ZbnssjbTfAHClEOXHb2onHF+4fHCGRm+kYJNw
BXkMlDRXjS9Vnp+AiMh6eQmcwQwYZ4curJkTnI6yr0h5EXHXtZAN0+l16QNL0SJI
9oSuEkomBXseSmy274Tzr9iobw0lUoO+ptKHXT1hDYN8xsg9azM7kGFExgfXr55j
dd/VjhI50Dx2bnDPRhjlKrODMGZycWu+ZtUSJN2WeXy9k5spdFZhzuuHxMILi4hd
o2tqta+i/On+WQ9a4EabvfB1en7Ym6NXe4L9v0TY97FZzI/+UuNiHGU8ldsfGMuu
r1Gb5zu5jfYLhqUjkr6azILHNnHL+RzWsRrPOykc4B7DPIUHZ53MBO7rqwytPh55
SmPfgyktF1YVjeK10isILL411EgYqQSuBW8VjAAJwl+WRsXsKR9TLALfdU2ApPWh
9YjT2BxdDklzCk7zNBhh5wbh/e/DzZ3SNQjhE8fcjyIcN8TOnhpbzJpP+70Vea/D
i6iSqzqbn92m8q26CNyQW7VP16+Naxv4o+CxgF5EADP8p+wD+DjQMsbM+0WfZZ3K
Knh2oq12JHrZQLCnynq3GEkb8EXPdklEtvuLNhRadlKgIDQF5thu+beLturb8jRK
i3kxRGIdBKlknMRB92x9YL/er5bHOTPUqYgeuY0rw9ETaVGzMenFAYvW8sNar+Vn
EmGz9ixX3JIu2iRw/Ic10SKUDJQKD5K531fRzdOQBIQ8rEKhluSAdK0PlecO5FlL
h8f0KdvtOEwKsqGp5P2jO1hACN2otsJ+QGJ/BVCpd+CFpHDhNNoT3eiI6Hu8Oku0
62+WRLgbI0b8SEIrM5r9oB3MCziBZk9olhUU8MnFYrNpIar07VfgwugauFOYipME
g/zkRrS1QrzpHskF/VhuGNNGSTykXHGP3BLWQzyT0uItxh9e4NpP2NX6UDgBZpfN
u6T4aWRffZ5yH05VFSAqyKxGJP+jpaRqY3lXPBeM/mL+mb924HlDNaN2htrXcBL4
v7sFmpv9dWkksXIYlfGTWEbA9qINk1bupIdLJannbCJAzD4pg7FANYd4oLtS2y+t
jVeNffwVgWEmXYMKF94eV31yDCQA6sldScj/kzKE7masuuuQtcFwGIohin0fxk2d
GBsL9tpjZ1FhoyCsL/0lxYP2wVdE2QPgLPep5edsFS7I4tq0r/WNhvPAif+BBWXT
TGzALcUJz5P4wHVBX4UJZxNh0YM2Ms+S5/xERYjxsqbNm0jTo64yjC72DfgYzzlg
NVM8knWfPKTiFNlwg0Nd2tfekr456pZulnA5oak4R9zluoKu4DVJMDP/sjLjuLIw
IA+nVc7hiFGYh7qM2nEwXf5Ppx5OrV2s3gsjSd+lM0FQxgUAwE9YyrpQNkOhCuTd
weuLSSsD8YER418vnBEsj8dxV4lHW0H7H9QEymfGc2yBPvxJW+F2QfHRw7F5XluH
ZKT5ljEIEghhE1Ilc9BMJzn4NOU880A+DzvfPEjbIpIdYICptI83ji9aHIqBDS8x
6CPXSybpUgZdpT+x6kvOi14OwcGx/L2UwqhxiHsMwm2ahPIcEBDmCsBvpI/pbMHL
V3xrrDoCrXaHe4XuTh7Ob0ujSUg586IcFRzvsNnMxBo+BOLt81OcgRHY+xS5O5dj
0hBLQOAfJAwkV0CSdiTk1GM2B+CmyO6NuZX12uuyptSESxqD76yfwMqC/HpvKKhS
k0nsVfxLrgXk+SBXY/GvEoGCk3VIUdFdd6txA46Taswm6Gpta1QxtSBoLgKifaUR
qXaUVWGwvTAQexYX6rB1TJ4I66FoqsH91SczvnvAKTHAOO9hy3E3+q75U8fW4qoh
uD5upRncMNfEom3KOqKjJ/rzlWIIk3dlqt/PXRGs3lDQ05UnxzeanzYILuBOwt4L
xurKNFc3vSYB2csNwMCkgFhMJhyQ61OCzumO2YzcXoPJOB+BLRvFLHr+ldmObfz5
sJjaCQeWRkJ8hrw8nU+n9kW3kYI1dVh9w/qmDWOnqvfx9MnrWjoqq2+RSGNmfW3K
lYRoq0VRt8X/tcv1neZeKJOMpeGKgEh14zF31MefvenAkbgZw4cZX1aThVGZB7i4
GxeMGzjfNNIwqqUQ6ih0J+bNrOO2xgz6WaTQ88sF/3Dfaj2VAkf2xjTsW14OPM6L
xu28zZqXiNh5IqF6TWBCHQpM6tdpbwedsf3vnX1kwTTH7KbO0LyQBL0aBUiN7ZTJ
Aoo4qFiqJf7HE9AEfKEws+s9u1x6L68wa1vXMsOwIphEz5MCqR+DtCCazkHhPTB0
n9WGi/EoEETjrNgCt4zd2ITdnIig5QCxZY+3qDikC8mvpcW9miqpIZDomIb0xzkm
Fnl2WvXVhOceOMZA8uR1H58Rcj0lZFQSavmrtFVy5LHDNuJnJRemFXrq1If1Hq/C
1WQLBpFtpvXF7i5WPWXfYo1mso/ENlOn2deEIXeXJJ/IqJtboYVFVujq1MrlMGQ/
lrriReprWrHDpmq7DLsGAO8L+ej/3qdt/PBO2xxaOiFfDEJy6Io4DHSzE6Gxme7P
DMIHbptRNhTd12F0XnJqLpqTd3/EEHEi8P2cgQ4vbDiJ1/TmXVMMaEHLoU+eMpG9
w/g5n/+3gzhAwO+4368cK0rNM/nQej79+/4MLtOia4oGAoExsMt9ibCZx1nzM+z/
te/T26HNQakFq8E9XJ2kTpGJDg9XRC6dbeWbZcsxN6lksR7s7R7rqsj+PESw5H2M
u6Zxarayf8vNRrxkXajl27LAnp7X8kFNCxZGzoemn51G1oxjCmHHoUbrhne4CKA8
8FEGTwkpKDnM9zwRsDYASdjisCSGbyQg5qIPEbM/F83XTuj4JA1d7Mrlpu+15dBd
WgBvzojvLKLlh1Aj4WBvKAmINbw+qWw88X9zFQuxcYLT/h4Cae8ORUVfJkCdpREu
eWuuZLnR0TXIlzOIOID51qTQ/3PXkDpvZ9P9zhpSABQKbfJuUtCE0kbJ+IMzdX+e
j5QRrMQZWcEXn8tbesPgZxy7L70YrKjN/mAnU1EjZC8x9s8EXoKsJ0kmp/EFi2j5
bbj28lGiP19cvueW34gZ5cl2LwEBXiqjcjSar+uniCs7POhuuKR0wMs11TqeZxYH
W3VzByApk5ssGus4/vRGKg1+MXf0kiT3n1Vk8MYbUc7gOVZe8ZXGl3NYmW9icMrQ
Ib27rhnYhh5socXg0pmVbOmYXhNIxP3nBpKkq65GxXceaQtFtY8hyVZHTGT4F7tr
FjiePPrM6s3/LmQVPXKDxtygBFuxqzs+MNGbeG3VyWb7OePjXoGtenoGNCWl009/
ZvawduzOVVRnBe7y0mIRSfihiYLB9qeD3hfCBO4Ok9VNjNVYMN+rjMIO+zVEHIn9
RMLjzSj0lPZMpGPcv670iWmX6PWdkIH938/+pLUtaUr2s4AbLuXJvrB7p9jU3plm
lvbRu7id6sezNGV4UIlIWUJz4Q4luqqNbiFnq0RxwrhlDdOqZsQ/dnlyIEsB8bQJ
Ap7NlQ6ahNjU+HYXHuq/OTZB0p6PUT5CfgFlaXDlk1t5Oeoi6YCp1S6xt6KMgNMt
V5j3k1pIXjd0NsmDhD2PU/mjHIGhMejkSEkUMsKdeEYL1lkUBKshNJP2og5hD9+H
2j2K5E9unmawonKV1WpR+9NYjBnoIivalZnsgncJlZBRZ5wT2oizKcnqfsVWG6OP
frd6fkbGqMw3W01Jh9D1QmB4v7pwvXn0RKeObyawvA7BAOtoPqQB5gOfWlzKyEEg
wVNW6h8hyi/ioNdjXr/dbtF9oFAU+KVzOvuCURQ//R0Kiau8v1VnMEgf1loqgEsP
XrkQ1EbfH89Fa8EfhuQrWN7ZyPICQoZQ1wJcmax9b+V8U+u4SMi6tIemBxKEcuG2
Zq9QCsQL8ZCqbn5g5QJ+keteN5JHQqB078JwgfWmbmhBoNiG4IttMU1E1arn4hox
EYTjPCE7TGzeAR6gkhSvoj+G8xALKhP+VFGlferFkPJHZNhGsF13r5f7FYeEugFp
xiu/mu2TithX8pV1u6qyiZpbIMLwev6wled5nhMfg1sIAEUkCaI3CqzDBeDOmoMg
sGmUXMoObuMDM/P1wejw3WaySnRknP4abC5YxUNJNDiE7e5qtyb9Q7uedKiI98Ly
0CanoNlh3Gj11tj6u5IG4fAHY6ySusGBXELS4PZ7WHOcLdktT3ctBc+EBoEys5w+
FOuAPMm+JrcEYzuBqwL1gCU6DKlgJXB7nbKV+sk6UwcypHLi6nAaW5eARwFm8gdb
3Uh6j/9n4g8+hDcWIdODhJ85VOdG9va9DQ3GOI2IZzbTzpTYdya9W9jOesywLYSW
/GsZ3vyOZPhsXATiuwhLyXD1aMYLlHAfoNbQI8FWgjqdLIY9V7XrmE2QjssTiVPo
xUEsffG9lQUPykK+9nYLUJi1stiP6hnAcRLDvgAsgn/+qaEs0Y0UD4VNnmRES2TQ
D8ZX1LQnpv9JWIXPS/aZ7Y1iz/5m/GIXdMwhYjaLaKyIusOQGMqj+hUdmpuFb/8h
vThjlXaVgaXtTlzvaIG6YsB2I62mO3UBzbChKMDZrr4WF86YFwXZoeLl8PmJAd0+
eOROnIo7uBtzibvMMQ4s9WMHwnn5qYLpVHZD+d+P5kVGcWxH6/zRmdQZED8vo1uA
ozDiMn/qzncCqBtdYC9DlhkFs7jc9bGy2Wok6Rfb+AwkNTkgFntW0hl/NLaBIQTO
Xt/8j3jGgAH4BwzB84wXCuZaW4tXJIWtzyDpi+VtWV9SfOhvNNBpTl4jbINMri/K
TvuMuPFRbzqDQEMnQtN9886gbqINy9OBPre+F/ziiPshuOkn0A1w2t2NveDxlk4i
UgAjBlggRHi13DmiNd2Vkb5osCRWlzsKNPs1my4gzj69WjDUCL3JxFbsoZBJ57xA
pDdmro4WOGi0PpHiooF94o5bQC2Wz0RATHa93d54CKq7wsLtXZGUYjb357+6Cpyp
zbXTlvOuEuvJ5GPFSYLRo6tlwKsEaKZTRV8bMe5PuESDcLO7i6pPF6ISiWu/4ICL
Pa4Cssy4t66IdzoXzp96tHRewa4z5VLI7T0G0WIfq3Fzfg8utUfVElVjAlUSzmNx
eLFMku3r5Mx3hwEurBe0CNliwQWXBATJbOUU3sHI2PWCt9/K+f2tAWXv1VOk9phq
3izBwDmztVM/1uB+h5LO3xc7jhGSgfvYRU2C7ptiQnHUVCCO5FLpRx5ErRyFVB57
AjsT8JQwMWxdAGh0kub9SSGcEz6cOMsFWOT5jSrSstdB0O5n6EyI6+pzNQwhe5Fw
Rp8jREtkVy4uYbUwz3B0jSMiucOf1u3bMbAuCBCSjZ5NhH87Au6Hbnw0U68TzJ1w
R6tz76esEX+VhcGFpYTld/lJY+9XqQM5M5bWEoEl4Hwhd8yP07YhiKytGH/Cmj/V
qZYqhJC3//I5ulABZXGV9yFn1RAuBdPsdgrY2D/Jb5u8JLPJXNONzNwUpO+Tr1v+
rM/YAdBH43Rzik2GPEH7gNYfWLxQuOYMSpYB2Ce3y3mn/1Ngz7VWm9BVd/Jf0X51
eqdgHxM/Z1at3NAovBJBLIVcScAIBrQmgYDNSbhJwSj7cRgDLD0Lok+9JBTCj5cT
n/mcUawbAKEt9aggBbLXbTwzJCnrMyI18eUJaPtoL56QcjJyGcCEugrpXi8jQ4ez
EFOov2ORMca01saC0r3bqVSwx6y8FA8bWgZML2tYxwhfwyIWSBfSDPDp1APOK79R
DjEn10g5ZKYXhxcKiLAKUU0Jf4JaAh+LvPIvLANVfCfail/5mxWPkl2BSmtEAIDE
QrHz72p03HtFTVB2ZvT0csrT/2H9ntOx4afvOliUFIrk3mGGxieIFKTGen5rMbgG
zsSCOR1EgWbYp8v98xoCw7y+Q4t1vQdRj7iGJi2b8yYEKQhfbotoZiDcSBlpwNLX
eDsLG3Vq1g/N102g/OLKDlKvEm466IxCOoxPhXNrQIbwi/WoLWZTxRr394tHG1hb
p7ouEMgg+1XVOmofQbcigDwG8Ft9lErf8UA3lGpuoqhSrhnPCbq+Oc2Eej+ldZ35
GspU6fXxmZLJJ3/SP7LuaV4NbJ7tBTgq2ufp3X/9ISM1Q7Or3yv1Xm8Odd0VqC8b
0Nb/fcA6G9k2/bOmhRphxGMOG88uMvbeDaBLfn3j4UqV0vRt6bndd9Q0kL2wT+0L
npGKt+R9xONyBtSHCjS0MmyaGO9R4kaf575rUPJq4/65U95HqRBHpBentraoseP8
hpq7PpOjVgSgjNnoV/9MOCFNf7SqLF3shQyWxqVCgetu3BilmaTxLvZ+pGWGjL6T
B0NE5+Wi2GRfNIwOuq++4mQFqN2Pn47cu/PJEcLyvTu/OQDDC6bE0qzd6A98pFBy
lmpJKAVqulbT06dGsN731EzIQX/knYvJnHuRAlyPfJdWzU9sCtM/sWS/Vw8dlc5D
qpPyGjdf5fxHOfJOnX/Km/Y/M4gRd27hMWAFk2mw/FEm1hkBzH463BiDJWJ/qq/1
QfrkF8zke8bdOyZQIxpcN1mDgMl47N4/RNkZAivJwZTMgzyp83rE8zuap5rT0ktu
nhnAXPcXIZA5VKrAjy0UBsP3FjruDi5J1lV4G4ZfMO7GSiIi+qAEo6uOl6sQxSYB
Y32NQGpsLZJFXRr4Rm/Ck5sOuOSzueWvj5Pgwps/j0JrIAlltGEEDlk2tdSR58qC
8iIwixB2hCJ4iXmOSX4BEMH0Y8nOWqsiG2kMNzFYJWkCa4yGXDU6g6biNQcr/17A
MzT3xOANmda3IjHbWeTX7BXkHIRI7yOyZp9buONjE27eOLa9NYH+CSWTnsTbXrxm
OOvqj2634xE5wJZxj3ag0UI6/YpI3+k14jaI7lGO+ob2nWyFdhTZJDgCAr1l+4E/
WquaS+yuV28KKWEiz650sl/XzHmHjcl/x4vi1PZU6K1G0mlPgLlO/Rr+1lONIIH+
I8sXIE/98+mZPIxha7dl4v0GltoVEG6NbmgNvZQtK2ci1WWgnoCKmyIk5r4yUlxp
QF+gwg2zYVC+iqZ8gH6GzWIJXtrNEp8PAxcp22t8dFLbelJciiRZ4uBUM+Ap5Snc
Dhix9WzRahDEaklllyWvPeX3OCeR7m+M13CaoVBxycWhylG36b7FEY+5l7l0Z8Jq
xND1OIWuxkV8tOoKgEzUjfCWV1hWJjqyxVY2xORv00QsJ5UXzvcrngAnSYhfJMRm
R0ItZpQcxNB1DMtJRbQML79REPPhYdzWGFTFYepjLsxBIVg0vanERkf//A3Hgmu9
hsP8NrXJZNHFCQGhonk+IWU6KLm8aJ87w3/WYtPCBiRGtSGuN+vImoLN2jcH9Gq+
sxzJ1YFraKBPaSkgkmWAVGkA+Y3GyQwC3GwowqYVtpuc1T7ZQH973BVB/M7OitI8
InkYOVBwlbEJ4mNNJ6Cn/+xK89GBAJb13nypEORCRn6/cjWvu7KjCZjAmRfB4121
16HnpXBbkebcf8qOIOWQyv3n8oEGeL0DHrGxiN+CRECjJ7V2GlyTnahwnRlCoOu/
ifzkyZflfcS/L9y9iAxUGcyibPhx4pMcC30BiTUZM5TGXclINjQWEuTtAQHM3ahG
bRd7mXFEdOxOfA8pJGy8lndC5O5aviQ2YPbdVEjJAzm6K8/28LVhZOvYtxHBBqnh
/FxJyxseo7x4EwTgzs56zGuwHZStPDAFn8siykcA0gJ/KS6rm3jKUTd2/fx16F9j
ZHaixH2+SJfeyKb3h5TEhPZlgxFP2uIMCUhUxXjUQ/X3YJ8tnuFS2YVYCUGXsp20
mRHNcuikO76RJx2Dy8FlVJVqhFK2f/XuIcVMPiSyj3m13vOQoIjih1MAQM9izeEb
WyKQfkWf4MVDL4F+OU8tdJqAVrVokWrHOgYoMcSjSAWIZWbBy77q74o2NllUQ4JS
znOH09sTesvDfzgwbH3jsDnWiSI9UJuiBAvX3EnLsm0Xw3C3bOJLhdbrW/UK+s9w
2I9QxIfbalVDVLb5Ykd4tJg8oya16RH4w4z+lxbazUX9ohxxW/+LCRLsc5+RMC4J
ok9dR6eJWqPhywtG5KmOCYOkO4d7DaivHTESfR5EjJYcrZzO9tLxE58q631rpVuc
eXIt299gTNo5Gbtq7aMbAi+z98nlmqVtUA9pqZZUCxV82j0p5YexwEgIHQb4xxzX
37pB4cm2CEL8AqBhHCaBFL2UFEXGugPUynSOLdfq07dCxgcG3esGW4KDkcD72ed+
2sugOPQz7n+jwULPK+Km028uGHf6YBF0ktf+80Gs/RKP1AS737a6POc5LDyDXV0P
p7wuOA18VrXQns1Z2xGgc2j2K/T2o3xLIygJO6xxpmhYp+1OQ6pNonRGGDNWmPTe
QqvClSoKXoiSrkCfvCQg6zpgV9XNNRIKenePaBNxnosF+s7dxhYOINZu4uHQyWK4
m8NXgl1OAysozlho1doXedtEBhxDfk8xjcdbRbaqUsuk6OIbE9veUjQxKqy+bxiq
gLm5TOiCJSQ8Fs+WM2WRKW/8LQfEo0NJeZ6KuYEZ1D/8Q1vnYkd4BVq/UxeOw1tL
Rq4ijwncVa8nFYUahcuOyT0NbK4zJbZYcxeM3qFy25Pj1iGbfaOytOhLT6U3NiH5
yQvAlUswdq8J1uhvFE90IASD3wbFXWPcCoy8F+pLmZmxo8cAey6Eiog+ZYyxgRwY
UMLEkWX51t1j5XUFu4HxHLAoRCWAO4cQAOlBQfmENK5N2zvBMbJI2d4rZ1kdMbiv
i2pmuJ+BzJAzXuC9/Dy8ZrYJPR9vQllkvSCfW36iwKggxgMQ56KmU2KK/OWKKe76
gWPvj9B9oqvsZZ52RgbdxmxXWcC/E2hnmdF/sBCt2ev20lbeANhjdn83YieP+RWa
4e5JkAeGLrc5AtnWimzvVV8/Zjz1RKP2IowqGwSCIw9frodyWK8dLp+s5ouOdYcn
u7aWNe6Pj9koyeMX6BHexHMpy0Egh/6s2eVRJN4Ta611+l+Br7svVqusOhQWWXye
ytTHrwB+hlkzM44pcsn1ElTvYbqIhuFp7eTwZwIYLszAknQSPVZrG/MI+WcceQ6n
5bz39ynyRkc8aMx8p4iJXk3Gmx51Yyeh5w5uOHGpBLG28aBqXWtFn8r81Q2IEong
RcJFQuB5pnZRsr2xgsHcC73cj/5fYLI01fmq7251Op7R1hbXghnkYTl8UgOpLutC
ovptXeFSgaP5ZWtYxvz6LhezrQnnRu9nB2M9rO5JaVbiiQkyBEM3I+RAgcsq8lOg
Sn3aCapl1ozR2HN+Kkz/s7PVTACVkOsvxw3uvoxEgAUeQ62dejE1YkH5HzaQHPbu
l5T9N+9I2UxCa4jL79SP30m9uJE5JnT1umnC2mjy7LdMvgDKBUAzwe9rOgSRv65C
6Xr1Y/Xu8WI3d+znWwCKHy0cwsKRbLatAO4XYbNmqLGZTtv4wWXLH3GtRgab5ay8
KcHpq6dS0qEX+R47WGj2kFnRoNSCtQRUXvlZZG60fYytm9st8VOM57JZbUWGSaVo
yagZsyZ4dC66A4n2RWcKHp+BX70KQGjvRFNo+uCOzDFBtpHq3SlgKFYCSQMwxKdm
ofEsAkQdXWY644aCzAOdYIdyAid1/1MfDMK0lSyzBU2mMVxLPSrBG1ZzPCZG29ZH
94BTVnnvjrzw+rbE9xqjrAOlo7rdZVy2yifJZ9lgFowcnk7xdNpOjyC9LchKqdB0
JUqjkCJWNXhEWoY1Oy3oM02H9F8PZNoL1MU7opesuMZsP0+KANymgXNdlw5zRzJU
dDKl1FhH+xzLlW3TPef0ZEzpsfNgEeFKXi+dLOUvpZq5+EKO+8Td+WbcLjYzvayT
gDscE0aSa13PB9u60MpE/62m8vqWXByLMvfim+OfXATIUviqb3L/p1wUovIwDCzy
sOm3Cc3aBUp+NSgoInGENAQrypEaxYoJmXnpgNsuDVqZI4JJZmi5k90E8T0Er56w
Tmu1nqFqC+HFpcDFSNAiJ3lC2iCsSPE0soC3jg1wU4bCKMjlu56FNbccjzxNMLz8
rDV2qcHvSkQC1JDmPHhJcoqs0ZVoYFiNhnhIfQzBtdU2a31r71aey6TOL5RFjoge
7A6jh4OzZKl8w08WKLpoNotqIskuqpcch/QfvfLkGWj0dqDR6Ojk+Wm1i75ZIsL6
Se5Lv3bB/YlCOX22WJOox2oAhZJVuVc4Rybw9Nes+EolOvO/Po3FxeZYcxsyC1z3
ZtKLrCnXofPG3OEUKdEurKcos+uVLIlFP3yrZ9Rhi+BOgkOoKcLIPGzCcT42dCTR
IEy1wnMd/zw77RvEVt+pLVSgQNdDbkoVj8MEKzeTYiTfew4ASfSIq3RRWFyqnk74
M0+maiQZsBf2KvjDq0XUTmch/iLLq0tUsOdjXQkGH2Kbt1rYGmM0VBXjECrb3C2D
RLEFqleShb3o2rw2hATr8QibCI7WKnHeyh/ArhWBPj31rPlVkqiRQrHbOevPnmFM
F52RIyeknBqBALA9QT5hrCKtY69YhW6FPJfQxwK3BVz0Vys3Jd5l3psL/qhXSrG6
8Xpql4Gbd2EHFJgcsTWUHNsKLHIbz4+5hI1cIiUVzXV6oQ14aexcJvZmUjlSiTpR
DNwtkiZUq+8Kxm5noAUSL19XR2kNEPZF7XJkrz8dCrMRNmei0P86BUh6rZOsIaHS
8Gc+A0UmFaCcM1mGDaEVASoCozZYHAMTrAMyf9Z9Ro/SubHeeMQJ5x+TxmEwIWI+
SUoGe1GVJg7pb+j+d/1R/cSJyLN3N0+4LdFqd7AsrOVkZmsNV+DxVHdR/E0xsEID
F0Bwk6H6WyKrz1bZD/SCVBI4y4QmHJUwXcSG/9QU7MIJ2dTRmdLH/No5MxmoSL2M
/tyPyvC0rLMpTo7AhXEPzpIrqbbdbb2dKqphGv5oPM2nj2b83WY/ER6Q0ykP5wnW
pKvvEckQZ8Hcr3F0+7+oT4Ih9anE24atnmwJZNLBEJvJmMAkp4JjBPnOcMvgpM9w
ZKzqLYegVPRclxWFTBqMnjJGu9mJ5eFcIQrNm+huOPBl+vAnVrkbKhGfRnx///ix
sBxkqPSYbtqyfZnVGHemH3ufWwNFeXP0tIOYry2hzZPgI/N0sLktZuYAGVv/PXGb
LheJNHU+hlGMWgzuA/xVvsMa+dQ3mkhxQOiBQ6dr1tgdTCXCRCjLBqphYJiml7s5
zBW5LsW4L2anQKcueFskc7U+I8fJe465IttJesEZ9+WVlh0VHBF19o7QwzN5fQNH
iQ2Dgi/gn4VSZ7lod5Gbi+O9Un6yer9E8i9IB/EsAnziKLtAIdrMd8SPmsro06HW
Qo+arVuDs0ZUYtngRtE1A4/X41/se3oL56uC/geMaHortgxLkLBPJ2qVMZCM9cPx
9jbyD7DJ6kFMGvB17w6bj7EFv/D3X5ke6aui8yXCjSa3i6F07RBE/GsB1vYEN6HJ
kWag/GOMM6vrp21Zt+QqT/vBL9Mm3aYr/Fy7ZJFM9K6svwhm/Mhc5CXRratqpTEv
NdsrUjbz/zfHCn8oEApwupkwvowZnBW+P9hyGpgN4njUo2Q3RSSKFDEzZCpd9C31
U+/Xk6O6tH6iqL9etXIhO3oUTi56NAn6lApqVzIeub6HPClTBwfK98zyy7BtXmvw
Y5RoohlUPUrRdV9RjAI6vPtzW/9C1LtAjf5UatfrUQynhsmh4r57mCdxXjgoxIDO
m22jHbaimezIxOYBHEDdvEHJXXmgpZbALwzI7VecTIMNbu9jOIqvYDbzRPLUsK4o
dxJ1uMykF9MP9eQfcUFf8xTgUVrYVGOAUfirOD3MVUj6IqLMgX9oP00WuZnfJ8qN
q2LaY1oypIfSM+EQINa19KjthZ9eKQmYpW5NKiUCvqgF8W+pJgPqBnByR5SxSKUd
vPetDdoKe8GF8VrDRF0LYDlhMDRKmoIL2qAMEB/YZuHGGqOivfNVBaJjzrEqPJdu
RD6mPESluythJMkhgBlXG+FyQjFXkDBJjzWTi90G/R2gfFOXOoSImyTRwse1tKKH
5EGba+edJZpoOJaB+esw3A56gAleqxtRqaD9NETjLvqZrRyKOaAfJwGoB0UTp0u2
KY4UwDZVokUsevepCfSVC80d6NRIHZAQiyVITuKGUq5PfOUZoI74l+4TppaspkaB
UB02ci1vRVljNvgEZ+3E6Aa6oMt5L7uu6cYrUEIFnVs6+qN+MgU9+Hj8qsqWVUji
Sh/MMf4ZipKcBMijA3XN+sSbxfCC/bWpVSYcl0nLoIRrBwvL2kq0wHxzgwT2Btp8
TM+fXavdi2w49Cfa/j+yXOrcA3RCTD0TRfA9Ubq5VrJi1DOj9pgQeqgeLX1hGROJ
hqdMphsH7rg88XwJQO/38SbFNw9XsN1rrdSpGDicL5joa2hxmy7A18+5K6r7SU0c
QuFooO4YuUOqFckLv9mVsW2x7qEo6Mvsm7Yo5VqEZJ8gixABYFqaB6IVLxYjyBmD
vuwk9TqZC8YGnGL+8zMW4colnuQD+/gM2ROmF5Q5CJDHingR6Xi386/etMRxpjzB
hfYxJqYokZaEnN0Thxj6PEWg07IX9VmvBjxl7wO2Apl3wMh+NLc35tatov0RJop1
ygWBQwRmffzGmdzN+qZenGhFNxh7OhO64nYj69QqdeD5K9gYxyGuYtg1J3nVwzsJ
7CGn3r7S/91ecMARn8uZL1cPccofwTKE0ZwOGsprqf/I7/fLWaejzwwTTKS2vVjN
Z/ab1BjIBglvEOq21Y85fYuaXHCB5nDEyedpNcF8brnhdYADL5A514McXrvHVg2Q
iqK6iQlluoHzcGpoVzpCokJGlgmiN4Js4V9ULrdvopUJ7ENolAAz/zRwPtq+MFIA
UnDoaC4KOIk3BQ0D+QUR0gAsYiOCBqJSVeeex82Yz4mjpzeEJezHBBLWAOKCKrvl
9olRj+zm1L80XeahA1+3AgwdVJfB5mQ/KOakmqCxGL/HqkP15+9lGS5Vd7K6xYyi
sxL//Zjg6Cr0G5G938u2iMFvXs87i3UfxrKjsrPOJjhBuxBQ4MZ08nfnHkCfIcRQ
Wwx8EwDsIgztZZ/45FgADkp+wYJS8UWhk2NWxLwei+ir3pIfFNB3cKIuLWdMkmxb
cHS+lBQ134eAxZKy5ImZ9F01+JJ/kmrn5Spl0/aKeSVf2oIZZI58FNJWQTcpzc0k
Qm2hCUnom3hXLkHxf1Xy7HDW+sMbkdffiC1De/9IUPkJNbPyNmHd2qqD67jdyn05
eN5yfUR1d63nXh1EIbsusYDLu6btSbqfYjToALEXhPoLKa+qocErKFu8b4LpVCIJ
oTXc7wPult7nx4I8c1+nhQRHoi+3bjTqBqDzvOTM1QF7NFlclJVGSCwRg5iFterQ
zNG+TTNl/p3lJLxBoOFB3D+CS/x1M8hOUY4ZUxP3Tw0QbAeoAC6P3Vr7bf/qt+zi
uFQK48Enzr5k1aXgIo4BphKaVl3dDDMIpu7zatjfJICtsQE+A12ATXczaz5hxhaN
3KuTVhaPieBePwvXS4EZV0SNBidm7k3M+Y6/L6eFlDtdsWJ1kyy3zOu2XCbFJie0
HKPAi8vpUqL9qmE7AsTv+2/0T49aq8+iSP0dawH+x3jXBEbxAw4mZv6CuUKOVHn/
Rf+mW2DydWLYb0JjbjUNLYeJhbT+vflm07qIXHeQsR/tAYLISkQDnmBCmXwp9gOx
EK9WQhB97OETnwbL55PSQuiAmIZAFCX8zVvlySRqfneQLKZCaLNxONMiAu0DosJp
GKHCgLndqRCYWLzsJ2RaTTOQBPCSgj17BOg9czmSFO7HsyblZcbzFwhvQDkQVkBU
rg9r3RLPfVCfU3W8bYhUB+jX4NlQdJwvNNyGIQzGhEOMaXDDQaj0fhIRgn+CKwlK
f5Rwju9l/IHLuFiyZoj7auhSowtYoa+UZoMzNhrFpP2T5/wArN2hRaGHZ7ZZEI8d
glQNcu7DH2aen08RxFvd0QA5QyvxTrMtNCp2ldZdD/vBXw4DDrKjigiYrx1bhETI
x4s2ZkpKlfpHozE3fP05GeIx8CxPfdEwAvU/rzIXhAo0Mt3/5MScnfKEY9pKFF64
gRu++FbBQBp3LGvg/ohjnx547BL5YjK3qJuDRb5Qj3anCTi0vTyocURHXv9lUikk
g9hgFYcyh6/5W8IdSIjECj4PVMBoWsLhtXr14DAENNHSZxvfZ1E+3lJwLdfqWy8k
7nRZD/OBiv3hhC6HKfIKBjO/eGreLqM8sr/usOUEtNGEzJxs+nMJygG2FF6OuHk7
F3/NRmb0F7wfd6FHkvabi6Av9sIDNrWquOjnKxuy6IAfxl08f+/fMm2DuJ+z4cB/
JhRGtlqTlCak/LE86IKUsrJZ7Zt75ZyNavmpjFvvW4CNk+Ys6hIf0/ySo8hgaV0/
/Xs8rBSz+NrCMBADOYqRTnefyFjqqr+B9H9TfaAYDUc5WWJP60bjOX8LAqOUem8N
De02J4eqMGQNmr8c5eLvHAevwaNTPmbkhnN/m6KJVfKieriISq9N30FryEwD8etz
O6U2wnAd5JhLOokzMi47J/na441M4og+tomeQJ6k+DC+BmcHgFtIe8NlLxSS3R+b
ZcbaBzvS5KvIBj0L1k3JL6RlgoE8jJKxLxz/p/ms1Msz9oJvVZS/D7BPhj9uDiIZ
zUEmRLeh+8594nxN/gDNKkZFPRvCTicqUyfAPvq3c0MEH1o1POMe/dYGe8wsIouw
NY2lOP4jSTarkCVqifcpQf4NXF7gO7BvsOGLYhITfBBAbJmEmuxYVjjYP9nbzbrr
Gn0rb1Wg/wO/ycMNffpEGDWO2Lx66CKRb4L3bSQo5fKwLiBlg+QZtYBIBgRTOhLe
FUyLtPHFWHLZTcQ5zNGoKYS6yGxqhUa4VaLEqpRCD50wj83DfU/QSRulmdA7USkX
1pz0vvBJlrqZUnbRsxswtP8igsQ0bI3YX0lceHI+H6l2AEkpa3rqMrlA9NhDvONE
gVRblYt+gH1PY/PGQFzUDMWTXwqrsOhy6TQANmEXVViMRSVZn/eyiFc+YymlxTz/
QUfQYgZal4xnzP8OxGxBQClryYb24ekr0E0sef40EiYFAmb7yDUvMGY7UkVjY75S
DTfyLbQARu+2N9a2fCulIN5r9aDpqT9rZ924yz5QsD7cbaVpB2KebJsfZ0hLI8Dx
ZfFvJsBWs2VVB5EmsnXEfSggQyXWjiFz0AIB5QEqkdDlH8J9dawY4Ov7EGAyYZzR
oxeMsqfUFwgU6WyhdthuvSlD5LAqhmbJNTR/2TMjDneaiNvtYk16fzl+m6W0dTuW
r5/dVJpTD/8nfbx3EL7HxrAkM8A9koKMV2RRED8hWebp0HDU4mvCjklAGtMbgDhI
qwYYCQrfs+kf/7UsMzM0VCrtNcp9L/fTAIpp11CTz1DsVMjGmshW6xBS47Aaq+Vg
3whjZKXmt92D1OXVu/McMk6anzrz7+dDu9teEmWBpBWV2MIomw5zACcfLfpxFoI5
2Q+gEYPbVMjxEbxsPDINvVN3Eg3vufELaRcn4pgTht/66gpdWeulLVQ8/9NUnu50
BXeVBTfPtFAW/jwtS+h8tvlaNkykpTMTLuU72g4Jz9EA7dv/ZLnkoXhYxPOY3EJz
Ar6Zra94dQeGiObeMUcnPYRfEsjGY+wDcSNlCLANwI8WLG42+Rxmq2mVt25/LZSB
Qu5YnNURUrBnCKDx5G+Zvdrl5BK5o+feua+awFaxq9/x1q8fQKum6zaf8tbxgtYI
YVvkwmHjEbevZx4H++1TN7nMu1a4ok4YTTLNMQoQUYn1AWO+n8Zv+TdSCGFeexDN
QdBCmivrL0+iApQbb2Plch2A9r7f+Fcgh8jCeTrzwOTXeRhwibOAvXRgT01uog6Z
zlxqfowfJ3PbPaumhNZs2oVYm4mAHG3sxsPYOUk6iFsdo1aBDeuAlPhd2ukVwoBP
d9RIdwU08iYEPgmc9kkoc7JC/EAVfK1B0aFcK0owSsv7c/qOjRR1USmNNYJxTNS1
iYyO40eYDWvmjZpBtEvCHKDa+ystF0TaMwMX0wzwBEZeQANmndZA+2Ok0CscbPr5
HtKP4SzNS+StZLWAtO7hLk1I4NdLrbkBTL2jqtno+woUDvoDPH33PZbN1iZNweZb
qDIXuIUPqciz6fpRZeWpyjCR9JxQDKSW2KVAp8ORQlvEuCexJtEbngBKzNGJpCpC
vifDxone9aYR0AkixNK9tcZeeRtHaA6WfBIUOhISXDnH2M6n9tayeIqAGcZ8mEge
6hlSHgi2q4GEeZwyxFrO/nTGda4g07MFxaTIRUR3zVN0Lye8N3Np+8pv8V+qPDux
oN3N6lEpfoLXClc9UpBSnsYjCuivsFp2nOPKquSgU8gXE4/9XshG91l/RpSEypSS
q30awSuTYGOZoiYfmkEypZbvukU2xRpm0i4481j+FVCh+1jl7az+bd2pIdkH73dD
1GYgYglp9/Pph0dirPd+k+AIFH5II0CYZsBRxd5F7aqqldB+8qvER8hwTigUCPmO
yZeUs4XSswTebBY7uE2FMaUR7hjscJcOho1+ST8a1AZK59eY46zVESAVd3HbMTTE
kDaM4d8ytSK17baQ8qoieLX1UGYihXGu1HxXCz6299CzcRMWWjTxPqpYwyRwlm8t
rsJ8FiVj61CJIafXrD6ve7kUxCtinLsa5m/xn8TSlJpKMG2hOdxcuTfDhtxqBzal
w04gFBMD3lObD5JZk1vauAC5z2d7mqQz2Ub1cn8wqgyrunWfhM90ou+cbsOzW2UG
I0xslMoG7KeddA84O0JV3SEXMrT2SQyoeZvIecMgTjWBG+Xl6dazqtrB2ria/Zen
dichDxiPvFiVH6BepiJfxmSgPI98ReEA7mwnR2cmc3JUoktZYYaDOi2VPdlrPwNx
/vbT2b17xLgkOzDoZXzTnEpej7TmyaUjhG8+PYLuq3WLd+sZEDBJ8pen9KysdSAm
UzODNu1LNKAJLNhGSG2jZUcgfUno2d51BttXo49Wx/1RWH1prK7etV7lIEbFTtLo
uqpYKar+OitCMF8bc2B9M9Xj7WLOPErKy6cnEXFBvFeJSInS6xT9cOtuYVFYngAi
0k5DX1FFc9wuEKaK1I2Oa59f+mcI2DUGXUDDY4Al0Z/P+ec9Aptx+mwctZLGmtDW
SzvPrwwtqIWn9VihUFg4WqBycQZJ5QK8V5wupQ9pdBxBnamLQc/QB6BOfWI0GcX2
rMHBTwuWEyLdfSDa6cRp5V5O9CTtD6C7pdAJz6SsyxJLInTiyn/pVN5UEmRe0lmu
uor/wX81YDUesj6V6QYPEeJ5O1x/0ULWlKm3fgDm+p2/7pJ27Nc0LU5UNcNB+2eY
4BZgSBHr980puHCbMs77ozKiRWRDcbflolvqd42a0BMTwezZrbwHPO+4zd2y6BTp
UlSsqwn3m0RYxwXuG3tz82k96o424/ayuez7yU6uxVkbwn5V+dOITtUkAUftuWd2
F1eNquHyk28V01eWvDLizzDz8rmGUgQbQ5zyhqupwlJZAt10uMdnFpMVr9o0JYg9
qFlPbV7yzAHyC8O3efSUVTLBW8me/7opWAJgw7M4dlEB2tgl2eZn8oZa/4f16iO4
GK6efNQVvDwDuo1ySQZrFHll0Fq2uppfGJH9p8ZgD8gZ7yh07MX+JSyR607axqIo
S0y4B9vrbnfDCJ3pIHHdzwqt8c4ow7oQf1Wos7ONrxWBFxb8QArGcZP2HeYdcENK
eon7YAWGnZoYRYipj9CztDNE96zna/Hi3l+/LJ/GPzExTjPY8dyE8nZy72pl8kJE
EGBMDBijGycUBxn/CnqQpQLZ+zY5ldsTwLEIzXZKr1s5OWBUUEkNoH/8gdp43Hn7
flTOGv/GZRD+IxFr53h6BDQl8abCLVeMMYq/8RKL7ebaY1ER5VdpJykpgYXSUNAv
zNI5EaLVxy1xZIEwxoKzslkqU3sKBCi6GkDA3CGIE9Ye1NRvvbrO5N3zMMfo/aEL
qm/HZZlqXJ/OvvdkdSUPAOkwn1Vs6+JXGp07MM/zukwYs06ZCegFK1zBU8pUke90
qm1y4yjPDJ14t0Uk5VJKbyvPvPcHfD4iqj2KACeK7IebcJ0HT6PQmQBcMdBPW3pl
9U7DNYf0Rt5dl00lDtZBxkrVTh5PALTbEaUGQYo1sNY6VmuiAfHMTr98bpBXCEGx
3W/yOTcKjTs5Fo3QTb3BFFLqV56hRvvxIP7r92SCfR1xtyDoUoRccNR6DLzX+SNv
tIh8LS+yOhbgjOjTOSls6E1LuzwMotPV7fkd9n+4gnpQpuDd1qI43+rFa3ZWoy43
c3NDlQDAn6pHM5BOKJGIb9kRV9PC/a8XfHRGb3bsJWyf8vfH/Eo9Xv/pTvW8obtw
s9fFwaj5lhFh8vutYyGVr+LJwfP8yvZATeZZr16tGSnVIvvEFlp1c7QURfqM62bu
Ht3eGa7EwVbK/bojjgX7lShEYjohq/RsfC0eoWxP8LrQ6Qr+s5w0kOS7KKm5jHGv
I0VEYiCx4A3mcOx8sMbpdnRiJecfOx7iRmHdHV6qAJMQVHXC9ZqM4eqtgc9tSPVg
mJX1hYn54FC4zu0+duWOmXOyKRtDA5RFNcG6s/dcRGYJQfVvWL5VyBvlqq7Ff+dA
dR0O8BQ+5x3IPhJ9JMsxpONTkOGSyAqn/nQ26H3z18Y448c67QdfGZwamBXpE4bE
d/kWEwlFUYU7knKdY6uQb6ihhnYoIF3l2OcC9jwFb7mkziwKKEVCVAAuXQUxyS5O
vkHGaK+pey6FPcYevqRQRv7y3h4nxSkaNngLhlI2OR5g6a9uRffr758A0rCTfpqX
+MEGuLXbwJ+S2P1qPx/pP3pHYXjYNskhxAYFA/H/xN1RAFs+PtpkNh5dWGVSCuTz
a9jVG2dB+gZSHIUYp4LxvaNGLpdd+vHw+DKqzOHfudQHSTHbm6Z77NLnOw4tce4g
7ndqaNxD5Sn1+7jwwXOx9KgMoBlscpjc6tXfjRl/QHLnXZHN+JeQH5tTzN34/dsY
S0rJej24IQXIzPIXY3if6Rx7tQaERq1ub0BEUsf4l+lhSVTBzXu4vvtjeA/BnuUB
rTx/YVMNne7bY8BFnUErFkiyifZRzMgbRKYpWqjM9fD7/F5u087UC2OJ4XdfJjGv
fNM+gz8uwZBRm81leaYiSg7NpARJohGbh5082KMexQtygmfgCzYR1MpgisnAcdVA
9NGPJFJ/3NpMggOoh89EpIDtrI3gY7ro7++uGpbyfG9ZoJCp1Gm/jqrfP7X2/Yx0
XBIeGkI5JNOTmTTmwfu8I3ueC6cLSRYtqNoXtFnILtDtFYVDRPciGm4molvNJEbE
pxdDPeXc7zxhylGH03AwPv5I/eI7zzbxtn9CmdspeVtLgsSiKewKYUrKIcpH/qLE
H8B6EMi5HVsB4fmh+1kxwL8JAjHj/TW5G2WTYftuuulvH5AGhVVPZ54PNvO1S5QI
dTrYuhiiGvLQ0CO9VZH1ZCH6bp7+yEsY/Tt37KUjj+G78hWad1qUdh2vY0jBu4WS
yPwze+ZG7AO7/YYhovY7IDWjQV40YhmTdctPieUzUUtwHTWgQ9ZDmmUsOs4Gyt7T
uS3xZ4kHNLbUUNKHtr/1w3Kanhbr1Yt7KPsZA0m7MvWQhEKFqA4OzuNneJkVEJ8U
x9TR6U7ufn1KupPrwrmnfO7EZ7NBYis1uyu04F2AGlE5pjiF6ajSYkVm4fiLntgN
nPOhQMLc+sh4oxYbSB0SCtopCoj0ua8U15ltnlDyGqfc4+ZlfZP5hPkFFlpBgiIe
P6XoQ8BJoGlIUPgUAiIEz6DQAWdn2CvQdIZYP1duhQmYqFY0fOCKhT4iFdxP7ZOZ
fCoihgv9/ALPZ6yj3qnkBj0UG0ydaLQ3KWEU+icvF3OizS1VsJowZ4kzLNLniMe4
CEsMeb3DtQAne7YvrI8mUV7Ic/K+MYXBnoTP+Vz9r/1JoW6NC+zlbC8vpGp0GiCf
FyOwF9th4wfoZ7pEMbfr+DYWFB4Cgpep5ZMKEwLYtnBdJBKHqpj1qwArgnAsuSYK
9bHQrf+ssU0sBFtnypTRBDkrqUM9SfCIa8K6Y7t4SgZO5MxXGbjXHC7GuFYuvwPV
dpGWm07Dy5xfOi7ubUEX6G5wKcSCORYmI2XTiCdcPrwtcdZeqrE/BoprC0ttjtRb
4Odzf7ATh5sybY9JdtkyZOfkVraI4Z8KhjuiF4huj317A0TNuUHg+/VKnL+KSyOZ
lELYwqsOTMN6/e271eNtWCQ318HV+USceUBJFnEYVV0qmOO9u6JaSClI/K2nfNxX
tYIKfkQosJYrwCcAsF/q7rTg6+KAiMvB51yWEg8OIuerKibs7tVk0uKshtB0BWz7
TdK8psdUKlZbKt9p0kFW/W7LYC3wZaeZSLVrQa5W/MF9K4bzAGya/IasnvAgj+cI
/orDVwB07xeU0gX9MMooh/jESuTfo0sHeUbFeMV3KyihF9QePS9KJWYZD4QCX18w
uNilz9N1n50m3miLDVrn6VKnZWvRTdB/F+vIIzSoBFQAh3L/A2gbV3yB28c6cLEj
gYdgSgvIgsI4BC3Cc8xlk1UZXMoH9X3kysh+Ddx9BSmScO2PbhTpFmQPRkomOPfV
Q7oJppcXo6ADb6MrT9nUJYPZTRFo3Dqejyi17SlMxO4CZpphAo7mP/zT/LppNZm6
GA5zvdlASH+EyoYnUj40+IZsFPWa8br8Qqi0sqgwSVQTkjPbDNUcSXtAnlS0sVEy
o7j/S1QTRjlBBX/WSs86jb3z2UgxtTmR0mbONOAzkmCgrFqkXcnbmjp3t7L8VLy+
q73JPMxSVGGlXf9V6oIpHkVvgn+/RDuY2z6JcyJEcpoqQU73GfpTVuQ8+yASn9Ps
gIeeeMvARgvXMB8mutluwQenfp3lh0h7HReXl5hI+EV/1nbrzUONgQ1uoIhp4pje
A3WPvKBEtohYRSOc2feWFZW5f8z7LBXcLIc2lEC7509FIX20nUnbQ6gaqE74tzoE
15FtXRvE8w1papEuCWtxo4dFd1gIhqFMPeQoxhn5HmSTgJSGxi0BkiwedrgO7hdl
tP9vHqP8Z2n0s20X1+OSktosb/b4VQvWVEeXGxuWFsd40kv1O+ZoNUiRYAFSsimp
OGWZ+evVaT+hee8DkwNCQAAGSBPrPXFSt+1gX0Fx4cROImLVlviUgMlOQrS/oU7u
KAzHZv/nw8PJ7vaf0QvtTTbrN9kMkj/Ye/vJZN1xEPTe5KAPnB81nOzs0YeSv7nI
yh/1OeY7ZncIGPh2TJRRtk0+AgegbTaETI/0y8hn1AZL9MBcSGqNQMGE078n3X2v
ds4Vv2WZaXGEXEfT9UntmhFzk9nSMFQ5FAfKCpF0gZO7tHHXbNluQz9oU3YweNCE
2/Qde53fcE9R52B+MBjmjzk9VlbX1XaXNhnlYXO3BHQkOAX71KjnITfAybxOcKXf
Zp7717jS1T01l8PefHu5KJuXTPohVHRIKE0UBL6paUV3VUHh9R+dGRr0dCB49b5h
ucJiD0+RmBNq2BNBXFqna9Rdk6lLVe6EgEONIeEXUD6PX7jYURBWd4VckS3Zlyem
ScM7mpQzdoH4AKDTXipNCcgfE9OfozyVwoSWOiRX2rMh/nF7VMIr80d3+iNf7Y2W
RNahJWnLQmkoGNx2SPcKXHkQe/lZKqkSyGbvND9pt70IgmuAr977+O6cFiYKl1Nk
82lFrVcpHZF0NCd1/wXTUKxM6yMwWsv/vv2mMJDcMyJFcO30w88Ksng4oao3SQTy
xLVqwIS/gJ9IsX3LGxhmyt4y7cX8vUniPO7TUFdp4UJ/WdUquHt0qv4XUjwmDbK0
vz1sKavBAJ8ovr/62W8fC6F1JA6i4huTzaKhsZJ9vx3uV29p059nWWzXw124AVkq
QIwNMDsv7J5M/8ZOLjya0vssDX0vU4k49JevD9A1YvNC4ILFthUtkSJjKXk1ooOy
Ofb+/SHTnEuc/fcLm8dA6qIZtts2nGlG4G9JtyDpa8vJUlFSJeZqNUgjzQ6fd23a
em7Lwh7TRB2VPg0RAYH59nOU1SJIBhkzFYnjGONba0G+LMfFdPFKhW319TSgZZyE
pPRpLmRpy3Yi4hsUCIikuT6YXjBdm0RtxVbyMyEK9Pg5rY00GKFRWoeVehyQxh5W
7mlaXzM68j6oHEdLTX5DTaSk8w7FTYUDHD9fv9mthRgoJ10smFYrAo6ECnAsSdwg
DLQmI5x68RQj+kyVZ7ycv/muDDTqnSqdi001THW5/tsWX2SOByNOiweTQmNs3kZU
4j0jHSzqyQCg5/1TXwfandu5ZzfVjncYyoaEZBNQRhDbRdia/lqm2g3O0yRNwER+
pN28Gi7MB40BKyrPVLuO7EO/DBtsWoV59Ly+awHH8H1fI/hhWkKBbkC/Py4eUIB6
GWnq4PlEv43Mq+SAhRQC7kPKgnctOZcTuIWcLPVQwJMJgfY5qZf1LcdkAcecA7Uq
efP1OxCRDMbf9Ps2OtpXhSazn57dQqOIDpw4p27sAoEVPmhpBylTKKt3+X0HTLtX
aZLTO+e4NdGeuFKFxFeyE+buOj+14YMzP0vQEsKISu06Dz22PH+qjtfNI+5Aa/hn
/XEq7JNRl68gubvlAkC42w02OIzNRI4IsTQP8+F82JQq4ea6cc83F1wMX426VsE3
+6rRZzPLjS3Ctc+sAt8ejjejLhBfVZ/gNEodylYtr9pLNSy1jk9fSedGUdYu0AQZ
TA8Mac+XO1HZ2Ypum00LJRLT06dAKTgFHF7LEx8RMNqGY0JB9jbMR06LFG0cP/CV
xtNVKcWjHtkM9kG4XROMwU0jx8zJ9J2piMqf6D3gO/gcovkX26PizSIBZpuL3hT/
xv2nALqr8yHy8+vzz90M0ghDlfeFMXAkcuTK+MYgYiLrKeRKNuTwKXCnljtLlKqv
ajVcgLaC4JrfHQ7Yk9rfS5+/y0KK6xhdhYv/AsLKi9uev3vu56KYKw0deOQKDLT+
7K4dVKTOv/DAvN1mtZNR824tEYgNuZCkKJ6Bqr2TCSnlc7XLDNmdXho/4bFL5RDp
5o1GJKRVBzhgWlbQi82Ca9vWV9JAalUhfKkNxRD62dNi1PLHex7yQ1PcEa3Fdgeu
EPEbDaJZbYtXvaBFNXso0ooyYpI9FF3lnEx4H0CynGLv2W1ZonRtdZhQAZpQK8OH
eNMFYcdPhzOeRVtg4IboWVPUrKqd+3Eryry/8CnBCtyHHKiskcoPDTJO+XcjRdrS
2MsT/O4emrJnlVqIhPfCwi4rtLxhvZD2tht7PYxs4szis9F00WXShgjkQJLJ36si
7TZyGt3SnQInwn5PmsU36e414z3U75iGmvFbwHhYJcHgLAN7vq1SHry6nOwdDssZ
KzZsPyOXnbklJ5v+trcbaCYwK3tp1/kMkhMy6wsYwTdlq3YMFbYiMw+/CngUnr2h
GHeUE4h01ZdnloXbVJVUFAZjw5kkIkayyMEH7wCqxy8qDc9UcMgbTkdJb29hRLUm
iCiFK/CiBJniNl0+mvLHqyjnWOAs0KpnNKU4g1QUYQB167rGvMvO1PAJ6gAaGsZv
Ob8rpdzaKGwQxfksfm9z4HCizmKNumV4Zpr6Wl5SBpQYDC5YWP7+wZ7tbK0U6n88
a3rn1ZZYU6XLxLm0q0zWjs/WZBw9F4mM4APf8ZUzVa24wrmBt3IlFcECxyhCmHh8
WeKYt65Ws6DrtaJLJ6Ex51XXvTd1QGENDYTsrsw4pgvKWoc8xDJC2ra2/9yvGgFz
L5HBhIGlhjosFQosHzG59LZskYS3pxYckG3leORmhQJKYPShl7AKYqBMLYPG1JhE
h/zRT2pouItx1BxoTeVVSPV3XBzwNRC1pwtZOGJacJVXlz4NtSAzVF2GHhRNzXtO
NGYK0HbMW1BO9U0gzcf7X/jNYiz3Ar88kla+i/6KT9+fKqBNgAcklEO8DhazoysK
d5pLUb0Mg2SOJVLkYCRb9bHP+OCHApDGInvqJgrOuOU+K5lvIAB5UGX8LeShh1om
IRvpLLBor0lG8+mwGNcdTNrVpQAkytWuRmetnCYpbwfqqaJHd5YBWZL4+AJdX6Fe
ZgibKqJaB4Oq6dgZLASGT21df0DHBfGqCQmopqNZtFAzLJxJTSzQlCZffKEFLw5p
DsdUlq7+t9hRFrbJ26uu9RMcEq9YXxFp0FBsKdQROE33l+oU4czNXVSUTKTlhhH5
9VpnDQnOTCNqBjmmX+0OebDQEFka+6QKHTA96al3BaW/oB8hLffDeA1ZzUgFgKx0
QK85YLC7Zwm0RMIoOcX9roj39mq3RWztZE6eiuycLaWhUiJGav0KT/oyU9xDVxwe
R4a1JPJ2FI8OjJlOdjWmWqir8LhrMk0d0W/i6FTiWwcJDNB52zHUVUPCALt30uQ4
Y4Ff3uBDWSXr+KemJqjM84vNmGO4ZvIOvsndZA/6ZnhogK7jHECx80UhCK6uJiZ6
EjVUgVZbKzwJUIndUd2VMaCtv503TEo5YB0faY8b7/ZV+QKnHh4dLTJwZcfMFqWv
duiB6o3mvsYzD/+CMJdAPAO4VO+JPdWD7O4vekKHf4tMD1xgPjAHHovDdAUVO7TG
mitRP5jyznlQNKfU33rZq+2qI44LIdEfPxQmlcvAiY+NKNlsbDVH/WYSmo9n+/Nj
67fGkjUa3JXp5nC84xBKX3/ndVqV5+j+JqXwjGNqIc+vAynieL3EVwzpzdPGU8iq
4cpAGVFHvbxLAWd+fYUCIRmgxG8wgD/C52oHwuKlEQ4EGh8CTW7PY8n+82P/g/9Q
6Md4f5VPz9pzFSyY37D/wyge9qoZfNPIkTpAotycESH2f+DdWgVcAuM90EA+Q6NE
OOnP7m39nDzLE4ulOHfyzCGv+DD4nd9QHubQvLLdqmSckr2ijT3/Kas5nDAegNNU
F4w+bEts/MijMbyGUrAZtpdjz6OljsM/QNfnLhqzCwARLin0PgKTDJHWf1vq22n0
7zhKPueVAG9vACjyJQm91rbS4MLRKIoAqptPwG8QeF4EEdFG6OLYoiVCy54hGnUJ
lRgyCuX3gO6B0G5dO94uo3qP0hIbPPFdR5t1C0u5IrVE4YtnVKrPvfxOpA1mkk0Q
brfG/gKfpYrozMdAg/iaW1KIE9ZIvpiJF9lZqpfW9kPxCCarBJS3JjniulwXFFly
7FdMaxXiejjMNLg78G5pIWxYkIuUaVF+MlCTmssxQlr4SU4qODkm89PHL6+QnLJo
kw2m+ZN3G//wjBwZx9iP5jCSh3DkBJpQVSJNe1jeFaJ3d/P1/FSm4fV8C+vb3I+e
MI+8gG6idGma+aPayCQRYD1Y5wurgJVQF2zorwZ1Wwn3abNEa5aiqWIekWduhnW/
a0uENi90Apax0ouwRs+fQ+HjT0ErA8rGhoPWZOxITyIneamFpJlaVYTk07zz22tq
taOgX/ghz+sWVyI3a+AAJ7El0K/uE0DJ3roYuYokrQ8+2Ejxxyp2Dk1Eow0qZReO
oLolIHPeYX3naVgI5GeswvnF9GfpSH7ZEa3ZgnNm/D0AumTxkB9Ly19+yf6QOAn8
ckRo82YqAilacS1OMxCm8P73qjbNJ8uRGklD+Sa/XAweIOB4UUk7TGs/mNRytHLu
fY9TiyEzwIgupJqAF8VNDewglUCHarIoTgJ3z4kk9dJQAgSTZb3OKsPw2oEftV6E
ZXtXvdLWWv7GTf1FdmIxkj/6hG502RUzMJDK7ccxzJLGTViEubSonpHqw0urHQ/n
bfwPX45QNqsCYHVE9cp2oguXKckgexzVPHeP89j6VqkorbeT4dnMfycjMdqMWqwd
K2Cr/h0SOkNDhz9EB4I5YptKrRXRWzK6R58iGgdip7u/sG+OCEkci/gi8xjk+FKS
JhRm6qqwHsNTjF6SHQYQ0+BqYT74RSVWKBnpZWf70Pp3nLexBv91RajhnY54plb7
eHCLG7WB4qJPdRDsWuRSDIHIUbjUPhRrAUkJTBHxhzyupK1xFckbUiucVlZbbi/7
9qVjPTBzuNwEFm0piJYKSJ5AWccYoCWSCc/3TT0sImHmK1HMGEVS3RCaAbiuX/EO
tD0Ds5O5gCPc5eD6H9C79RsH/lSVsMcX3ivEpyaKBY4c4I5wl8t8gKirOsZmVcCj
HKM83eJYeG2p0tV9nEhdxvZ2lZ8eTMfsm11WiQupyxGrUO7E8OQj8xNmDLqWqtP3
EdO5PI2/c6ps5tF82Trg684rUyQpJVWZKTW1L/aXHYxPyDz2qrI6L4E0ksyUe5zw
ZFSc0gO0GPqN0mOOV0A8SxLV1iQDOtVW/M40qCb5HUYqR0gKwGcp9OkdhmGNKzkE
YcNn7b2er/+8HtZQkPuFSa7rgwGprP7NMCuUh2k3eP3tKf9LBBm6w8pa2KTw+I5q
Phrjw0D6j5q/v5td9NWSNMO1goIeX3r+1scIGMaokZX87P1ymyoX30oZDVSBFRpF
4abENRw37FXQDQJTdADSkgUeQkvTDjRM4EXZSJZQBisVmGScuJj2+JVbaXdZlOMS
QUCYnjQnI7MluToS68s4oB8UBiEhz09KwM/YjUYE5LAp5nwNMZI7ekuCgzOGka/5
0sIM8lzITE8F/K78NF9o6bZyBe33+6rtI8y5FiXhPNZKH3CqZLVKrpeY+nUw1GMJ
P67HzWjDDZ/W+pvipiyfuP84CHLHhyFJfKuYsPo6ulV+Y2GZ6rXPL0wGLApwJMVi
5lOQHaScJhnWwga9mBMyi+NKWP7H4tYJzJohSKolJafVKy9bLVX/PIsH8dw08rbg
jxkUl6yOuvrLM9pxLNdjJFtCsPSwwsHWRMxB22+GqXQQgvwRYEfeGkuwFTuwZRmS
Ip9mOXGKAzcctZ8bvXuP3zj/6TXPtHjuW+NtCz/M80/aSGptYLCB0KxU8+kO20u5
0vs3DrBhjlr4jNYSVLHTmKpZ+Rj2TSOBfhgCPrX9x0Bt0r8Iv9p1cmKkNHHqXcqI
Z7OoT4Cp/u6aMkCqQTvXI32s6hSIybE4elWXkCmeDlv4rht0swifxYouY2vPW8fe
RwX4ENCPs7tR++EPszWKNNOox/iWl9KE8+pSkE0AfXc4TD3Khd4tC5wV1d1fKq5y
obQfL3knB5tHZ7FkQh+5s+5NEPmoLt5pwmOn1mLe51C1QG2NvuKsdzH2bWPrNK2u
x/eKTF1HcMOYUkdfRHxsfapHjHXB9XXBRxevLezZcJjoSS8hIqmTatmzdMDshqH0
6jBRSKU/aoR6VrzmhIT4GPxwy8j3WXN61jGrBy/0LuZUCA3JrPozzKi1OpdLqNXS
dGBL1iM4xb48R476VGp1GuRItY/TIsY0SO7McWmOjNCmmVngqBcpMvOIgnrI0j1o
mvxJU3mkBFUW0kvrusdBa4fWNJHUltvUtgAj0lf9kkVhPa118dyPx90BGckD7HNU
D7rKaa2lsvONAhhh9S6ilerYL8n6LIPbzT8NuwtBo9i77dcEB5I0pLPS6gxy3mRq
akI/NcxiUpnwNNqmLcuN3lK4nK40rItqBnkVI1S+P21nvDQ6Dtm67c4lYzUAuNWW
aw2KJxAfsjBDsSDLJkEbn3zP9KTLa1z5dsxfKIJ+tsRUDqFrdpTqwbfz6+hiY71s
c7NoeJvG48a2Semyv3wIktHV1lWxvqPN6BgV+6K7bMVQyYITVb3iv8xcuA4f+AU/
+KKNax3dQU3aXcohNL33n3q9wzzYZVerjc/lAUPYK0IwlrGKl8N9YQrBo5SZw/vV
s+agf8rXFlYFGOLj5KL/Je50TZXjH2VNoAXRbFuqRFIkKNrLILY1JlUIZM8zZprj
C6JuXI2QZHtMyqPE5TbLd3hkDs/Ns+PoBqGQF5OoR0fcHUpQHlPUm1lSm4Wf+2e0
QFBkF7ZyCoFHCcFYU9JvJE2u/0n33rLSYLmGFBY2R9SfZSJS8HZs0xASeNuJxS7D
MMtome6vr2mLsdZjPpJrsBEhPNebSaUetqIc/GrGH+fDeSkXUGtKKqbBrVCagPjF
gN6N/8vk8wcJWMlXzzglibmrcuOUDmTC+BKVYlz66n1NWNBqFfNzL2U/BpTjn4bo
FjlJtX/+pgR/St0JrMRkaILyXBFm0dmPtpwei/+kELt8IKnh14SwdDkHA4JSWEyQ
bqMKwI0UYfdUO4CdRjo9Q+ZM0YCSnBnUEaGIk1vTcwccJcBafLHRbffXHWkZE+IO
Hx9UPXg2SsFLlCVXn7KGGCSCFxN3lUgHgSsuDfIcJeAxN6II3bA/6YDs4lD19fbF
zBbshS+uYSpiMzZ2n9jK1kcWqRlATxaxA1VBXQM7knz811ecX2hknQqaUeHyQ2sE
X4TcJ35QEXt0vlLEQVaXvRQsQoAiEv5S2BoM3HYmmZxu5rnXv0+pt4wSgaN5Rfs+
cHQIF7iwzxk9bf/Fm+ITdKcYhfQyhGoB1UOIvmyJ/21IJofFfwU7y8ClDAsRGiBa
BbQvXYR3/guSdUekB8fVpnumEutlXi/8U//vT40u0g4rqfPDbQaTL2VY85UNYCAf
Oj7TqmJmUgP5FW7SIZY7xmmYjHH9WPtO/RPYX9IiEgJaKqFwjN3ePQMOa1heU82M
od3SmITTgY243RbuvjozNYL7f1lUMXC0G3KsHCJ0cM+37tRutmlzF+awxMLPss8f
2hmpKZ3yjeiNOr4EwxeKhxSFoKVfEzv211j4UuglKqTlUBVEyX2A9lEP19/CCkwJ
7KJ8Vu3o+YUT7JS6q0LTqVHDZi1O8ySiV+wtoLnT2o5qNVEQq1O+2xU7ORCllOTG
7x4+D1iXuk0RVanwQv0TV17ZEIf8qvlaNcY9yQ0uaqH7MHrauFvzW/3pTXItFrUa
dtj1PK+7Dn141nNfCQ5EzfEFc36iPpOG1Vgr6Sj90yE3mvh/lmGgyNVZT4doFSjk
ld3dqrLhcjOtJfP7PNC69vr3qPkU1XWAVskXSuaevzRipXWMTl909frPWr9Jj09s
zqXWWjxR0E8OdPyNB1AC6o2u2xP3ZUFZuhizsThDRh3Judg5idx7gpiPkDkp6TpX
sXOB8r3YF55gBVcdav4scJLDzYNI8tws+VJTXhbY1tFhP7pFJt4frLa5SmINj2ZB
6pFKwKAIOw0zqqahPieRAOTCjLQ2fGpo1hVTQzNJ6EnvF/U8bqunyyLVVBQ0hmow
YgEjllZTn/05wOi1mMpObyOorAjlhGjIbYkOVPIlV0lMJKko15sAi8LEoGCVcbGh
/k4SNWnPT4Tc/NTiSSsJedy4BrxjHXajbTaA6/uczDtP5/J9MRY1Ze9GVJdVq/6r
5KD2TXQDem30/2kvtW+sPDHMC+o7PG3Q4pR0DGkYeT1X9hw4W6eoKpUvxQE1AROH
FcI2/9BpfAOf0uejcWJVqbkx6BApLgobaksi/f7H5nxFrgGqMFq98TT0YUndjYoc
i+eDPw107RH//PM4vkf3FwOf9BVjVTLkMMrtuhHV1we2aJzYclZ8Yw0UJilmq/gU
HQ7AXHFsoog1hy6NHTxg/zPBYmEIepc1OtB0SBfA1d1fp0ZF6TXrLh5JBwjGOt71
WvMVBoxNL5fx1Ez2B2iR43Pu5UD0BF/F3LXZXOoWYk4H7CGx9LlTXlBN7YFaj5rs
mORawfS+Lf8b23V56aF0xgkebC3KouaRCGeugH3oJb9MgvJ3E7FfjtxxAvp3kVEU
jFgDtxONta9aJC/6iP0i3MR5ElhD5oXfkZVFGk9GD7j2PgvTYa+yV+yPFBJxDvrp
sNoH13VU8TQyMdTPe1SrRXD46wLIuPap6am27pSIS/JJruLEqlihm/838EJjGsmi
0YF07Lc8dVlzPpffMvO52q4eXr0ZHVsHVIt0xE/+F/L06Yp3iR37VmScY79JhL/l
HcXFhT6vEV/LyzwLqAQGaSTvcAJW6svQoJTP0kr2bMRIwtH0/xS3696nOF/9i7T9
y+elD0uOa46x5UscIDmodgVd7x2ujmc2uioZi3DwbUVa4/mCbj53Sst6Nxo1Kvso
b4nieFcMrwHYqxbYxZ0q2n9cXvLi/FjPy8CLFk3vgESjySeZwlqE7fyy5ucmntW3
TUXMJwFbpLjizwIZJtIV6dMZoBs/pJ3HeaARKG8ZVmQi/h0XqwWOdv+VPS345iKz
ctjJBSMKeGSPtjOCBbBgny+v7VBTqt89cL8JMy2v94h84ss0hPvQ2iqQxko+TEzb
A441gOkhfzqWWQGHAMkPqUaU613MgTqFaAkbeLmdBejZRhGG/1X/fGSb/yo4NYYz
NRm7uArCNfvFwXCzMbaC4oQvW9g9+0TQWLY9Pka43pol8tJyai3Ngp7XIds26/Wz
bYtxqIm4L5N/WGtNgHdRdWzcfddwtqp9RQOgUkcF93GgbF0fnpnnzApbQKqi8i9J
61YD6a5BLRv6tqAt1jJISwWwPxArqRSRzwk3CaRVMHra6lvv3AtRtr90G68OoXXp
JnHgC6Bb4JEtGDRFqoErfjixJgwt1LaTZWYWx3gZc2Q8PvlN+u5q+f500FWxGBOO
db0piUCq7gVGFL8CPnvUgzmXLkPkzs/DFaaufaneHTlTWRrNoY+dZRnyLlyx0ARa
g8h7YF293WNr6rvG4XIBejCe2goHG/MmOMzKpWWMRnzLFGJCgnQdz59IWD+dIGW/
3CFzlWkJ4jUqJYkfqbQBzMHQhLK6SH2KRcvYoXdEyVc41mREfe24mKY22XraCoF2
HEXSigx0g1fAe3M/rP7qksR39gG3zNVcVPh90SFgQBT5HV131ECg7ebksalDmXmL
vswG16WRlOtb3sEA55UruuHEdqPG82Q7dutayJ6aPzCncJtrRtNN5YlmbrdIi9Wl
BEyTYUJ4zgxcEfP8wdPh/DCKc1h9zVQuSdN3TVK1lCPsUYXDj9+BVBcnC5aqNkqs
cfpePhpzpSiWpv/+2V2QbGRbfrW1sjNBF83GT+1mbecsu61aQuAn/A/GCYRW733E
4jamsuEYaePCIBuEhKVpDa/yIWjpSEmRRnT3nZUo/Vbl4i5h+X92PznLYkIgCCQC
U4Ts/37zkEZBI7pqcX1V3sY1SnO3oKYDKIx3MREOHsEIYuERh1XLIyfN0tIAceU8
gdbzsW4nHcWw6+IkdzXB5MU/tBHJcCF3I/17lWloLgmrQgm1faABei4MY7ZBqVHs
k6B4TdQ1WrE8SQCULo6g5/G9SbIarlGACcP9xF/3NvT2g9noWVbxHUu2oYxoPdjk
AvKonm1PzjT+w7wZDybSE9sBc4YZiB2difKyyUPsskLBqPa5HZFwGOOt/8kZhB97
+moRxehPas8mCFBNx6pwIo1Vi4ZCQokIlnowYAdbHGuzQYaEZcm074AUxqGoUVyE
1Kcb9CILFImnNF1fxuTIsVbQE7XtkRK6Yjjx8WThPn2d80PECHEhP3tbPHIoHbgC
Cx9cGVe4Ha//x5TDPmNDffDoKKzJpDJE1kvgTDARYIFBFb1ZG1XZrazK7570X8A5
RGfKhsHC3vniRm3D+zHErlicRoinB5e+wH7c746LndRBrbp8xk7u3EnbX1k+akqX
de9F2i3Xu/Zt3gavZoFfkAtsFnGa6zkjlHqZpcxDRwpc730ATXSpZED9GW1rna5J
Rr5W+5Mfjdt+kqAc0kPXnF8IAKUlrc2qZoP6cMBtawj4+B7Mpq4Y+CoOwC3k0hzV
VLrU2sZRqKdoJ1C41TpBPmyFbx/YHia2tmczKZO3V3M8nrnaImsrgC2QNzQrpmkN
Udl5Eu0n9F3Yc23RPIxkzu+V4ai+iSApdOK8HbNtt6wjziw3cK06xMEvaPhVZgm1
kiUYDNlOqesC1/MpmDLYvajkiNz+Xr7UvVs87wImYo0zZq/momDE7kUCvltmlX5I
JI11VOZsUBZda89AoFdEcpfIL0dBtRt4IQn4OT0/Rk6xsbHOLp1Z+lfyV9ssot3t
D+R1a1lafOnfe5mz5UPEdx7GUdlur1LGd6O8KfiGRYiikWTBmnEaoWR7G2c7RHxl
yRADk0DMmnBouCMN/wlXuBCeeEIBi56pu4IDFok0YiDjSOJbmteyvlkvmV77dPM7
ZFor5kC0Ewv0RVmSqvzmTYVHFjnTcjQmEu1adPI39AxUeGm5Hs3iUhX703gy0TES
VJCMyfS/zvF3p+LzkMvYltunM7DSUK9wVFNzy4GEjNhb27D0LMUaL1XUfuXo/gn0
gjhaV3LMcmHfLiP32zPfLf911t7PH1DdzgHwSRoRuDFIMJO7KVqelG89MpM9PJ4G
HyQFgRNPTbBo1wyU8M04a7fesbIf/YWBiaaKTVwfgU/t/dx/n6FCBXKsOLEQpZVV
vlNgDlAPE/w+rOV2NlkhrXdN1CKIIe+OsHutNfy1NL1jRdWWlG4iifGlOFtn9H5Q
OCF4xICr/Wz8eVt00HfP6lWsQ7BWvyOOcfEfo2Z5/h43wPrFHLTcAHGi392AWXU0
lbxnkkL7Q3I+lzOYFugB4fMAo3GknvdYW/KGdZ/CHbmEPiDV1r1hqu0VQsuq5mKs
Glh5xbdsif7BKusgGOgTjmXkxxkI+9tZUa23Beap+geV936N8DKFmhrddZ39Q7AV
lelTqde07gPnws+4lB5wVkIGht9oPJfHeWiKnee8iZVyzQ69Uk+VB01q/Q3MdjGg
GVU23JB+Q/yS/vmyVZwzDNH4xoO3WZhrYtKWv0atEIRQoxzrFem9jJQIhC0WMxNS
MIpqWR8iqTvd99nYFBkUOfJAmwJez+nPRZs0W5BH346mlUbPZaynf3QCsXWjE02A
5Thhsc9p4uTrdVtvbDG84DDCgM69Jb5K6cY9Fx5wSnfr+2B/N3OI0d9LufYN1sb4
Lpuwm+Q6yuemQV2yiRSDbsCmxSe/OaOvJtZEwjTHbE/NkICZg99ZHhAV4bLnaTI4
1f8f7U+6IuX6U7qLh+5UEAn3AW/p3SUpgG6tixGnKQ70VBSXYGHaiW9UYVF2gjHh
tlN9eKYLEJxnQ9BdK9BZ4O8Z6R+5FYJTpe9VWihQIsI5wGLurcyfs9UzuA1KxLlx
h3VpP3GPXjNkkPwbaCQzCG3ywE0jLoAMO6YASadZALFNQdd+aYdMW/7thth0AIZO
p9D4TcD/FkYdXdZRuBof2DMVDYTKWn6yoRuYvjC3G2Jecc3yRNfTkjKRnwF115qW
VzxuHml6a5cjnNBDy5KFNmxocHG1SO6dXbpYVqL5NzklKXI59udZ9YM99mS7dE2d
jcr+U5+ngS6k2B7QP+J+0XmtCPTnBaS7lj7O8lZLDFuSHBEvQxj+7cyxKYLE4fgz
+P+zxGAg5WUW6F8ySgfMxeYCedMm7MBLBIOqY+G/iSCFxraP5Yzf8v74S5wtR9dU
30fzDVP7Q/rzQT1l+dcjIZcVBRuLODuHIUd6VufFv+qruoiKQmdjwz5TcOj/7c4l
b7wigDB5+aXiyO5Yv0O9+lkSEN6r6OtsbsWGf+H8hvBMCODaaXofpwUzVbXSAkK/
agTobIuGmhXzNqDyBEFFJG9hrU55mGoeWl6cYBcD6MYz+oqyWPLZ7aQsD1wMnp/e
EHV0A3E8gjeTjCzNEJACox6Lowhl3Tyq7K0qvLpUPcFJou3FSLmiAmwbl5HuICue
NgKGJJ3dxRzqMkuiF3/tASFuMCvkBxwdLCyJBXuzzahwiUBxgg3rV44KuuSq63Ho
Cz+j28sG4CEoe+pGCcQ5u0a/NnoS9bcXRxpLex8i730CCbUPMURA2kpqV/jAM+ta
oF5ipDEnm8E0TJ6NQk+n9ZpHB5NrWWT4ZDIQvhPeunNtbZUDNZZMBh98Up0O6exi
VAJvnrsRVouzjrzImWDFe1xAz9ulPhYYg7sBv5ioigkZ/SureBbwt7N+kjltWBdF
DPll2iHk6EnQitbmHKDogoSMBo76JQxSertGawvzZJypDZ/ezSjn8NBB64sgWsNw
yAIaX+EuQQeSyhmyL3yZd0ePG0Z6HxTcT6fVfLh+CMwKo4baj1fQnhNYxqO8K/Wb
ABQJh+Gy+z6gc8PqB6E8HbwXxwe7wBh4/2o3sB3HRn823rNIOaUdx1DXQyxUQE9v
7YEXaDKGuWaeMHCgifaC6s8EiVBvdktko6/CcRZvWhOjG4F3qP2A0OJsXeJk4szr
UbcMWG/YaqlnAcFuBtxHDt0J+xSoW5egbp5gr8rzPu2bTrqx4jDk79+/1XEjREGb
BELJJvUhK1Kn5KdzVcXh2P4d0WbVDQ/FAeTiDrsw/jzorLqw79tYmyl17fIO86ya
RimqZ+YFlvMlzk7zdqDbLsO8CFuGbb2ZbLE/50soKkf1/Nv+kZKprZ/2Sm4stE4r
et6NSWXzEifJ2Y97nL2c+MZC1BpMFkwVF0w6TQCN6x39bj2rZVK9F1EEKFASzNQR
SQ/3E0OYJfo9qOwwRsWyVbir2JT3tuX774xymObvwakbCYJ+APIxpRj4KiRf0htx
JuqYyP2wm93C0ILzozpiR9cT6o56cRSpf79QS8frmAUkK34H4mHuiBEw/bq0ux0B
i3f29ShBuQ3CMSdAo6rhsAYSzjxnNg3rsxGgZC9EOYx2aAGGHKf+YG1K7wndhloB
LbZ4ePGAcAeAcnTaKI5D76K9lkD6/0KqLgmRdQfoCuzxm3jXSdHpN86/BmEuiBk3
kp/gooaD0Yr8SZosrjgFMTUAMlqbX+ZRIqT3TgH0xXKmU4VbKzZ9WBcWR/ca2Cwt
YeltmD+t7DWP3Cj5XbVwxfe2JhlqXuxWlFF4C2gLCIITSUlXinGIEv5qx0I7wPCM
dK65q6N78Myg+GCMy+oxgEedfdsVEnLvERuYppZ+kYlYNSbX7PlTusBf8OsjF5Lk
gUd8ht7mG2ZI6EOjreEXIacktEtjR8uT3csiku//7H6DxziFhm6S0GpDYbkRZmIr
DUQiCzaD2586y2y/Mv+VctUgGdx+m1OdUl+/eSGIUd2ulskFv+8/y+/LVo3RcTzH
1d0GWpeAsemwLpahzHQfoklhBQ2UsFITGWMTFTUx5ZByQ+aaVKRdqQAbUuxCLmPY
CbkoUHW+lTfOQ4UZ8gJwoqyR4ifLSyU7s/y0Frh8nxVwjMvyGmyDfcSu2aigtAr6
3lWa5VAiuzRUhSar+f3MBr2o4ff40772SdrKCmB703+ppCDw+S/WgpIJ8piY+mxT
3/pCA4bJprmeHzDk1h/qM9pYfxPnTlYs0mgGpgQaNdIYvB1a6HeNL7ze83i82Eyb
oE0hZYKpWWDj33bHEZ/AFRj+IaeOO2reak9ZaINONp52i9MOepluaeTQYWC784tS
wOJ7raGH+1EVoCNo9f6t5qqxzbfC3i53m3flaGeStr4HzjuZDjV98jB3Rtu2ozAM
jX2NjKt0WQtKlxYwW4F0sIngYg0UNYgu2fi35+jgA7sSEqquff+ie049op2NXPgm
zyG4z4giv0rcs1Zd1lO1v3j/WcjT2rzBzBCNHqgC/TeGNklYHuAK9cTwtSq/9/OH
THgd0WGhjvl3LqzbHVSxu2Fc5xG+AQqMxER4kuIE2g4kABAIfy+i4Ya/lWZ2XVgh
AuTMwmhQ96L7u8DuYvZCc4QXdXt4/084pCbwP1ldDQ8sCDvhvdZziTP6KH/L5GXc
TC3hZGKuse6eXTasnkFk+AxlJV0B0vIwX4fXEZFsDMu38oy3DG3TT3zFnbPVqlxG
oxhqNnDqkH1LyX5X3bleAYpDnNbBg7lgANMtSuAVLvLVAhncSJFL2fOjdQNRFrOD
gL4t+5791aXppofbs9h65O7o8WrfQ5wrs6YNho8QZB93sX48YGEe/oItxVJ2YZot
8pa/LLiPXKbwceK7vTjYqdwsTo3MFpd8aK3gmsCoh2DumxuKqqoUiF/nB+lRg40Z
+012O4Ygt5a7FxFeFz3qLajOnCJZ9fdOwU2NZvwLCxfIPNk2InknoXpM//1Im6Ln
3YjHoT0Rk9Q9OXMZxLXB/pbPldM55MLerix2Dp8U7tZOgqPfAyX+92pZMy5xM0Kr
J6PifSOVov1oiwInH+umtj0Rll7q1kjG9VsYDP88FxJxmu4d0tBKMlrT1QCVvW7z
uovYvr19rd7ZOMCzw1xBG8/OX5b+rh2hC/h90tI+cc9a8FA+Wml4Bt2EIIRYYUeM
XKlkJ+q6pJK6v0Kjhz2S9qciZKgnisVf92LXFFk4SOCKWnddEXJckpdaSwHSqjNm
7s8IicYY8C0ir9Q+4DvnXi/CXHF8cO7VzZqFo6a573Jz6fFDbdMBg1dfXta2Y7hs
n6ZID1av1nx4jkxyriPPp5hfFrGUVStahnVM0/mcEbTARGUh4E9G/w2QwLuBFW4v
5e1vFsOhDN6jFN2kzqEOltvv7nHdSkH7tRoYqS2Tmmfaz0b6OTV58vtTlMAFsn3M
e4wsOWQqN2CUAvKwPzVbAO7M62ubqEuCxlEBYMRmckEHI0wPjo9Qm8Cu9kqxEsgT
WYItxm1F4MI/8FQS0M6jV0fDPvovaxTUUL1HRrEJkvmJTS+H5qkv4n7G8uQh2cFC
jcTS9kqnrRLqvnSNTlvJUowFYFqStpWT/L5Jg4WGM15KNtju5gAcIrKHCM8Tasn/
49PQDaVnqg90hnpQEoa5SO3I1rjLhJf6PaOAYr6idu/Apofd8pyO6deiSJWFg6a4
dZGYRRVHQaJwc9ATrZ7djKEYfjn4kbnzq/wKH9ZYP/6nw8GR/2uTfuPSsj3dBoce
mt2seOjLnwJI8jYAXfkPhUcoZXTnDOKGoYkJihJyYA3zRgXpoiZASthz6fMgDFTL
VzixwL4Z3WhRZna29m2HAx5E36s1zSRH9Xl/V6NRLg2fDwoFuLYuBPuYXhrxmb3/
KmlFFtkLb1f8XbyjvryIcjtDECyDZDCraJjMDVHYq/qDNJbLyRNA1EfLtOubFp6L
Iz+IM2eqt87x3W4vbiuwJRDFNpbc8QTPzHG0obqncn/27lLBMQj1P9Hy8FTKl6SK
TIMp2fnNcTUoCUBG9j1qTIXc4MBBMpTMrP/MOzEt6tB7xrTHUIeJ1q0LfS5LG64+
ysWxusxN1koBlcL8gTN0hvN1rd2IlZm861UmfozrWl8M/Zi2ZoYaM3ZiajZlt5/N
7L11I8STNND3VOqXvZKKA7tWYQJTUxnSMJm4y8Dx1uU8I6KCXmnRLJJoVTLx+IyS
VU1Wq70sLNEhj8yC1gYcSd5G4cLIEK1oI9KjJOmgcgBTzPgaq4UO6xoPOulkxilt
wH+Z5G99UXxbb2cCbNZXnSQTkV1xXopWhpcMVhLHj4nNbpqv8aECdsu0CDMO/uoG
er8eyCdeLdTDNtgo9SZ2YKTKVjTKGAy1SJVmDU8AiouEF8SWoZaka29T9UjcxHHZ
jilQMj+AK+2SMkOvgAZsqXNiP6LisF1hmdJEZ+JuXRUalDcbXd3gS7jj+K/d9h0l
EuGrVDRsh+lSkh87YMS0wmO0tJ9p1GkfP3IU7pMd/ohow2b+kE111YrGpj6K5Rdx
hqgwdpE/Evw2SwiRO3QFqwugcFFNoLDUjbxTJlT2aHS2w9zTmS38Wsu/R2ba3KBn
+ZOD5GHJfiwYAHAXRiEfoJML5b50EJv0UEQWet7s4d+eGt7dw3IIa1imPOITz1tO
d028FunfuNQUcb9hprodzEOZxQ9lCaivNp4L/QASAyhU7IYrG3e2Y3xcY7KaPasK
YBO72kCyHVZ6jED9Ie+TkoNq7hlgO7E39IbXfQ852AeU70qtMLbKyHHIZMuEDERf
pRo5YkjtWrk5fIj5lx/StPwBuUm49dlIxilkWrO/11zTpyRS4sCXKLRFQmD0NeZF
AhArjow13PBNVOigEZPo/LPRMW46NgCnZT61FRKBFz8OctvdW5TjwnrVOCzxKIMg
Olj9VccTI9bIUXpaO/8CxdzFRkPb01ZDVkQ8nP6HNBVfhNCm2Mip5IHqtJUbAeNY
pCiqrQ+WyLIX3DJHbepc+AapOWnPQztEV9C287q5hxaxJ6+KNKYH2vhLfjZeC/Yx
ur5PNkLWXgnpuNL/ul3WZErt9uaiUeaRGvWsVE5VHWPYyY/TSeCXdtq3VKL6kGFi
NZlS2x8BVSLPvYcndhDU5TLs/IpImlfnxDPc/cBn1ppO0qHPvfMJQzpMOJSZM6oB
jB4RndLPqB28sIZyuXrolnlCMfyWziNIryJHIdYSeRYsXBeRbGl51sDMMBFJbLpo
bJo+N7w5o0iUGsKLIt3yhg9Ma0m+D3enegqnrRuAXNrF30CtnrhLpFNTChWvJu0A
iLDBKXtXZX9rAOfBvaASpEPVTOCYwKOwGN1/sveuhD4S9WwqoP8pY67fXgHhUYBV
/RBwlG6oMnU13TlLBbUisLk+6xzzhNLl/aliT8zMnYOb09yqM9ATEgY05CppWJpc
kPJ4qTdp48tprTgDImhPflrhNmBWq0ICEku8UJQWp9Gn3hATdclrcFcAQAQlkYmY
ePmUMrKSFDPm+x/0O8R6ZLaQvWJwi0QI+9gdDdqcI+IpwWOU8U5eILQ7t7cp5+V1
IWgJejHA0jbsRyRbv2I89EESF+4Rd06h6czLee8gUDp0OdTXcFQ3VgrbirvBcj7d
zbCjeRwz6k242E+E0karzlQPGdiZrdoOQiL/UQU5EPcTARQF82ex7REO8MoHOBEW
10TRRkWHBKPqm9TOZVWYlmUWYPRJ1+INiQyDSvnKYNz7lrunzd8r1kXJdyKfZqG2
7KDbQfGNSID6IZEqHub8oBljV5p2Jd8FJIaApgncxjOQpAai6552ZNKiUTKtcpkY
jqLNQ97nNRFQtPL/jIdZMjrc/YB3KBHn7YrnEo/UITSCG4qQEQatZDMcVlGA6vgd
j2DCkheEExvoth6oZu05cUPBZ0M4IhdCSU18wZqYECS6nvzqFmtK+2jYVMwY3zly
EtefCo4YzWSqobY+B3MXkALjlfbq7oEBctl7YXH1PNeWRXSq36qqkGw1vHdv2LNU
8vcOtbyg7qtby5ca3sfAioA2PcqH7jHDYmxV5x7CTOOUjgF5QhBi2hIsrnM1VcY5
XNXvk3yFyoLtyF+656AI3OfBK0R+u1vnnPlC1k+N8Nru+BvXV6xYsHXP2b0KZTBb
hxG+kanNb7rbUT6vD2ZbTQJ5eimoqlSz/MtNb1JRCEI+XffvhXOJ82MlD+melt3B
9snxBw0lWji3xTXHNhkBvFikmLGcTOgLxgGOoSveKvAjIPVhlbsP+3cPGWdRPZue
ZqgmCJ958iAhhzlrJiO1Y5OM3L5wD1uHaGs5DZ8B2xFEGGhDh4J1ZMEHivf4hee1
BSCPJEgMZ0+aMmYOaoB71lrxsoUup+jK8Mqh6LJLfv5FSGZebKKiZx5XVMDO8Ji1
tPZJ7gd/chO8avu/x+ulhK2UXZ21EtkmnJn+U9bw9VKiIcaKgWNZLfiKSd0nJXvJ
8XB7aTWp1gEGqHfAeGjojvNsXDOUOlp6m6RR4MjeM9jm1rkICy00HL377rGeTFSd
8F1glsEwoeVfssY2Q4zh6bNHb3sT/mOZmn/mw9QZT0Ok/rqMMOaykKBGLvGnDWmR
GNnDS3BMfaaH3zpFGHy+xc04vL1k777gGiTKAKLX7Zrsz+qJLGl18y65T7Wezd37
aQcdPGjTz3qOQMHaZRQxp31Yisf20kEF3XmxZjMhopPBcH4cxCDaknjVZkhINkYb
dcjdA7sMRySEApP83XqS+pq2Wr885ZeA/32TucCBVjX4kl79DtTa6tL8LvDXyM5y
Z9SOe0rMsRF0gN4+CzILm8SYxGDls+RasCcwKboaXsZTbNE4oRIYRVkvPg23M9PU
Ke9GIANLAn35UjQOci3Cr+BKS+lF7Z+FnGfQ7SOvti4OdfMX5nW7Suu84GlKaF6y
sB3eSFfboJv7kG322rcV4cetJubxqbu69mBc5OYMMoTptWYPnJrTV5G54HPHsh3o
ZHY6xTtn2X+/CsoRzSnBVuL9l040fXOpMEAP/RMh8orU4U+s8ujaKckkRgDFPWvh
vG8TVlf2Yuioh7+czSjltIO2vqGKcy4dPIFexBORXmrbVeED9N8YP+CLPjZ48V+q
AJ/X8Du9alk35TH9BIHnY0BKswczR17oC+Sg0y0fTryK0eT5jmq1gkHQBfyb+qxh
skQf3PZjvMyJRc7D/Bdayr+i0HNxXyaIY6ixXM4ndo6gaGQyDQxYY/BJ3RDlapbL
bkmpHGF1k4X5FrmH9ROxQfEcHNXbF5jk7THgH5LmBSYXVg53zoG8YPWB28p32w2c
w7jU/ZUo0VS5lZphb2AUGYYzgDhvO+8qYXF78OW2BdTmfPlWFXDPE2shVTc1SUfj
4r3Va+rdxseGyH4FUtVgpvAFSiXihcaFU3sTSB0q5fCUdfiUEI3fYtNHbqI5HXF6
GnXQrMye2necmtZxGMteTzj9CXHvi0W1o6bOz3MiRXGT3evrIPS/wEwlQcVJ7/TG
XiZmMIsqbiNTk0r7RVn4cUP2ubRpG/wVe7SadVj9LVmXu8sOuC0mjfa4Fp0/ts+9
pWye1owbroh7fjfM0/TnkPgPLoGqe7Z0kY5wLhgqKvIMbTOVat3etMs3nscpvD2j
q+U5xYvNHR/MCXi3m+vqIZ+gkYpE6Yem8PB/OUjK1RE90saK914UZlxSoW00vl0K
Tp47iVRniyRYaAE0MrD0QycFzI444cspxQZnGv+lrY7LIHc/lf/dO2jYGObeIGwL
nsSB+AgW1dVY/hs/RRfO7nhENVBUpaAdG6lsEVF74lAKmXYyUIbeDfHMaNS8salc
eP6KQeQIbBMe+dB1oeVp6xlclQ6mJbAEo7Y+BWP9p0HHhme6HtsCJuhFrq0z/zkl
ua+DyzTEMXHMhKV15i+2+yKhnFPV1ATCMO3AlQ+ZwhPrTX/hECp07Zhl8U7dw2+/
w5ddcKgjUdCsavi3eLY1dYmVU1RShOkw2v6sb5Ne1RZ5jELpspeLp6LodNLiyKzK
kbAleo5/UabtzbSvb/fAwcLgrt4Eu9/hC8cqwutHOAxj4wgwr/kWv3oYAGgKm66Z
ltPt3lov6mrabn16hgQsutLk194BgNgmaUmYPfIngx39iwa2gII29hCl7iE6HUVO
F0hsmSmYh1psed9ZUtu3IWeBPOvQLl097/ISxBHyDivpRY1464L7njrZEoryn/Hs
J1QFP4nxzXJlJKiAX36N1ZPuPC9qkngkhe3f0aDPxVKiIwB93eC9p6LqCHNI0Oxe
kbZnmDLFn4nxmr3y9vt8Z9mllS+7022vEyFhgJsnws1VZ/HYEr+o2HSdKwonctvr
MfLniCwvjAmm1gL0puD3/sDo1KX+0QxVU1F9JCQOvWq+qvl4dn6F+4pQUryDlqM0
HSd+s7IgDGzCyZbRZckd1ywdzaNykkaCOFObxCs+7DW9ziUOB5RXkuzU4i6mm8il
PigQkUoRwdtkel5haHt27tr3DrquM4ZhP45R7YTuMKntzR1PgUUu/W50au7DQyJ6
kauqMoJBIqNQ0HPNvbaGJzk8padAbdxZqSX8wZlXZ7l4/zgz82q5VDSqsSEq1pIe
vFWH/Jy5JRaeIsiQdmdatq/I93WwLwF8Te1Pp53FPh17E1+AAe8zpeZcvvKVmM0u
wjxZwtDhQ28hygL8mWqwJqRpX9jsypTyCutiTbriqdDq3DOXbN2JItLvwhErO5DX
Fqr1pW4vLQxzc1nTdzL2h021DGwpYPVwHYwF9swtLUbkhRodamL5TFXgDMEPBvfs
ZnBB3sLaV+7vnmSTEm8P7cEOAKBJKuPWIfcNZqrjbkSRl4Lw86Of/DqyUsthZDEJ
1K7fVfe25+ZkwEjjz8Jkt8lQR8HzhcoKqPOy3/5Dh28UGxunYncTE4PXNniQruUq
p+xbkpnjW1Rqy4zkQyGL/EBCoWzQTKOOH6XQdH1GZ2uzbaKpKU5dlC1qasYgeod3
gBLlH7tPYqecxhZOZvjCdYKVMehGwAkCL9goaxtRfRXKPRAylRLH1Vj85tAxnfdC
xMkXW4I5xlULYRuj/LfwQ6aesdknRh72QpRMEIz5MnTr27b/SvJrDW81o0b9PJxG
mgpdnsCS0SG/oRnhf+TRoZp45QkFBxr8ZRK7f3+VuZ8RpdTKjs++LSWXn8kbXKns
6COxziPy5anuQwSHI977+jMgRleuat78GPIN9PT/2RffMhijwCNLFtz2cjMZmhtv
KJD82BDAoqfsCoIxNNI0KAJUMUrNSozSqUdI3lIIne283qDt10GTBePAyVE2K5oq
1m7nm6KjSyyXxW/fQT33SIEcIdBE/1OrEjF9RMfLD4mhzCPtfYHuRk1g78dfRMAq
gVh+BQ2d82M+cXsUoaGLjGYDbO+ia+q/ajdUMGzq7NG/hP3tgFwvtHUWfYGgWfsn
PGf/QB3vM5IiBV+BwtVUuOvB5sCu4tisz5Tl6+3GsnvMyQipakSN0XHWXK4O9e1S
K7BVFfqGqh+hj6RFn8OJEbdlv5VpfU1SfHuVPY/guXr5S1qdXrJvtTrIJI0L/ayt
MPPZGe6hYLn0wEJTUWOVnQQPhXrGa4mD8v7Te0DiInFRignNEsG0YIho35U9c1sG
mKwYCCALMvv4JMnQMlqMW+OoR1pSmJ830qQXkF+tXJdAFeSxyAiX+MJa/UJrqqa3
aLfan9uctzcgV/+9FNYUL65CKeT/T+/eyQwEAbueEixumleFNE0DOigUlwEu2Kzc
gXKrubYBKTodsdRFIypfZ7ZqohKV+wqNHHLJJk3Vn84ks8FwTJxUwYpbPHbQA3e3
+gTF823XMQ5ndViQlu8gKIpNwe9tpVXZ3pDQeOcZtK/vRAiCkYfun6LsI48OfkhA
GIFeanVSiH6GiiqDia23Nyv/QuP2/2F8i5yuHlR2kIfSy4GEVzvDQwEmeylRpqse
bx7QAFuuz06nZqsLPHvFl9kzSLDVdU4wKPOAvAHb3/PAJOyqvSC3oy69LJ2Bf+Yw
uS/+OjwBEu6H+8DYhSqfqLT4yN6BIa/1deAweNCtgrY6I4ObeVpoT09vCDGdCv7W
z3vHAVCAebHwWsqM/tDRDqX6tf/RQ5ks7orIdSWmf/XuKZkPav94UdUd2eX5suhm
7Dr5/MwX5AtIDL0pJLjZ/od10zY6X9A81+0D8+EcJebZtquBvbW1ni/rQ8aF3mnp
4sART6HXVlUwrvDAeLKuOPT65gGJ5sh2sZGB7mqAvpmXSyUvZ9z4ey1U1mMq4sDZ
cbAaaM0Z9MJJ8ebq2Zr2819jZGYRsPco/AXWQ2xw4oCHYi4o5KiquqwSoth0uAbQ
P8CeJDoslCKQ/GIlJ2wkIRkz+TKo8TEjtx9Wdio5TFspHrZEf7EdlWh+Wvt41Dvl
tZVzHbypBDtk23rF3mWM5ya8SiBmewi1oD0o52XCCsszZV00zK+id2wksGymHtAv
zpq/D/i76K+FdAHISwlgwt/6f1NH8JjMEdgU1Qilv6AnkF1C8jmrcdiIdmNUjZPS
qIp7DHtku+sJ9gwElLfP9ztt46cVXMR/4Qfr0234Q1Y7wzeR9DzONQ4AtmgurBe8
urTA4ACP022+nkbf/w3UwG01hgSg9tABPY6z0TE5rbquyiAJz5yojVMtR1o1zBCD
5/WMwfG65Os9fgZVmEtoXpusgAY6Cbtk1XiQf8/5D0PmIkndBDBeGk3iGC2nazT0
HUwjGXWvlSgpboyPPq8rPg2UNjSZtKjG8CpcmOIuIoouLcBdpyHmgiG3WHAgCugf
yRmxLPf9dldnJijii82cjh6h+LPhrCKRZFK3s5WuXjOj+QZJJ+ahBeaE2R+aTNP1
emDDY0J8sXXqiBeVjvuTsLke73SODFhM43nJ4w6yK3AMnlnmDQIwDrT7t1x80zsA
qIrjlKqsPlw0NktEbwfqdcyQuwh3mEQHFBqUtgdk4pcUNpVcyDt37sdcD4bpyl3o
uspJID76C5B0Jlek7XRkqYDNeekubsdeuXFAoEmjRNQ8dfu+qnVDjIjEIY+dZ184
Y1jpt6WxOLdLotBKnMTHNRVo0NulmyyWWTyS8jdQMeoP0QvXqbukdKnJKjlCWCrq
tBGjGQYLepRqVH6m41qtoR2XfItAKcy/SMPsx7wxav6rr2//oxbxF8fPfIAuI8q4
IVJyi/xgHNrzGlyWxxLxdDLQncN6FB8+2NvWpfa6EYYDDwl+ZJRdNPKVMYGpHCyr
v+ArK7BofDV0Ji5vSxz8ogUgd2aYMFGGj8HcUzevWtRtzA37G77e6l8y7M9zvy9T
4H4PPvdcry7Bvm3n5TZu5IUpkfQD/j6kj3bDDgVCaaHLgI8klezT6QL5sb344HcK
7fhV8BDk2C+F+JOireHU5efqWgAmTokyemROCdDWamRa9CqRUdQ+LlGDFMdryWZT
SB47cDn/IShwiLlbqXGzjshNXhmEgj9Yp/3UktIln3liIJpd7c7JSIuDmiDFK32/
1nO4oZ2HWgHFyxbHjLUj3G4DrbKDwSz4CO+wlXYsmkYFYnlXUMyZl83n98OSf8CE
1oxDWaoSEDRzszwZ7GsLAQdp8yip/H+JERFW38XfDmS0HGwMoT7yzPk6dqIodG+f
K1tmKmPOEzr97jSslD7jN/iA5tRP9YR4AVf5XnYiw8NWl0n22jBzcnj1lwT/kBcC
42j0imo6KPSBUYi/zqGh80yqgyfLM86dN+UXXjHLHy7d27asoc8fEfelA5PdaQKA
kT3pWoT7pnFPCzML4ad1QfVs9T+8+dwShEfQ6Y96Y4hMd39OJ6tAnczSf1viZRom
hU9trbr8tDZPSTRYswpZwH3EhOdkBOcPZR5vNrkTCoc03s//l18oP+vXfVzAP1n2
8oraxb01FYjt416aV4bIIAhD9BbQ3zm6jY1zSQJRrKRXVKBsq1US+DCdm9hZ83gF
O7Z3anwcQggbQA5aPsNZ//rClPZnhftQ98R0onhOWiq3AfZzDSBfF6pnAZDCByc1
MXRFqDwCfOUf9hm9+RMEhudjSAbbnNV6iOQtejxqFvMcjOrRzQ08xGl3rDRzNFp3
OfMMWfx6kUehjAZa8ZQaPN8UyFfaii96vliv+SdJMS6IQQyyrc4LsK1opuBmePFT
u0zEi6fddIHthClu/wJcX+WEib2cy3e63k1O4f904Fu1/a4JJY9pldWXVL577jp3
lUnYlCRvJ0p2Frab05mKg/jLGCuagFFCIC1YX3srrRxTuvzWSeLnNDCCr4/rDTSD
/mY/SRuyXOy1G+QDDJZLOcJ2QuXAqgdoOwrAYXQ5Q9LdQpilJgenhpymgV7mwUnL
jEU5ogKdZ0tVHzGz52FZIyOFjUN+KDMkgSykCkLWDdoQK2OLCiNhLFmL27y23q4Y
hreOJ2x009xi0qWvDVP8TOhS/p9nbFq8NZdzuPOMd1A/woSB9fyztG/KQ8lvRL5z
A1fkQQIQSbnFIzxmDHcu0arTXwZvv2haByJdOW3A0cnKaW8idJGb3JTghmJ8Mgdt
MRodDJAe7kWANardp3sqbFYOGNAuNlVr7HKf2SbgJ67pyaEsyRuVr+qhFEJ7lu34
veci8okjfyn1fZVm4l7sf7hkfFwqw7WsqB95ymgWgY5XlQ+8QFVsn/jx6y5M3xqk
DncpeLDxgLfT8o/KTiBnODpbWMbDfpOEkYFhqmzVJeyff7ILfsiJgM+Wh49sL0WD
+scUvlWuw9a1OiChS4W31GMx9454Zc5CfkuIXzRAH763kvVLgsGjfLwXRz65fjK1
7Xs+ykxfjYZAIkjR1dRRCrBg9mw+oIctayUc3gZuWQ9+6uYmBIrv+pz6Bkp+KebV
Bl2NAWHXhFwq7KgGH/DRGILr520HVEO+nnvcUVKVZk4+CaAmVjKGXoORr0+HjxTU
WOKRouKq6qSSWgUpWq40iHEpt5QAIRVouyhpo4GZPBgNO/VHwI1AwZo5kG1QaRs9
zXpCM53g1UXPMeVP+0w+BkimoQaGHiS72UF8pmD5ikEQlEOyohxj062xjoaxN8yK
vV/VA5SN6+JH4VpxobaLteeasqQJtaYTSw5W9ocHvV1MpiKeyR3W+HWISFg07P0Z
AFipLQDFCKvG3CT9z40Ob820jOmPoSZQffBo9FoVuIx1T3c8UxLDch5jF2kLaBi5
FHAegiz+ZVA3yO3ZyYjeZJhdwGpsC5whjlXXnyANnU+EZfooa/3hMWoJ+WTMtop+
0OxhraDSIQzJrg81wtkBJsJ4BxNTfYn+vu28+rLWahQ+TSMmd12aWeqPbEbZ0ktJ
gtTL3WBooVr6a+TiRtqAJPQd2CBGvd2gqpobnl9NUKsMHT+ye4sbX4qxpFJJu64q
z8K/JyKIcmEgkAdz/PbhT+sgz/tuABKzmsys1HcPP+tIpMN+rPIKKIXtIbzhSBsK
DghRupRfdP13+FlvRSd5/I0psdMSlI6DeJS066GX4EezzCl9nR5BoYZ6AfKZQ0cn
UkkUHwBUSKRV0T9mEbOs3GFKhRiqBDc/a0+a+d6nnfqdcwi4LLIbY9ABcAPcG2VI
5StRhZtkxuM71xGgM3CnJGpuMKv1xjkII4mhwQDlZj81wRi5h1MGKq2SlcwexS+K
Ul/HWmmrt3St0roQMpVOiqSzZbWpJfWipSoIvPip4YQ7x+vROqgbAUTZLsUFpXT/
aEj7i0Nr1kXo2n136TVbChnZxtxl4ZjRDVxCnK767rK+jA4W8EeJhcSBs78jVhB3
7lFyJk4/EgFaqQP0Bha9NVOZVfGXFeQv1AZfsGys8fuJEKL4O2rNtb7Mxg34JBOD
6rqnFg+1z3LP3aOwPSKHBRpedPTtjJQ4/7eLO0ds1AnOjq0idj2ppsaRoNeHzrvl
kylg/NiDurInwF/Lye4j5EVqozUi6wo48FZ89muswVqFNhFHatroUJkQSYIzBC0M
d1fnTw84JxPKsTLNVyrLUF7QecXLH/WyIjGwGDyk6tgNCRjY+EGfxiIvr2c4/Fd5
hT8yWqWwaHsO2Vy2Nd6k+C4A5eE388XnYpwoy0+61n+rmNYgsABlrNRv8qbIGXh9
hpUGSro22860gwNRMudVpAqJibLVTTfYs0jRjLz+sQ3N7No5J9UJd36vgDRt/2y+
CGhZiEy0UNX6i4Vkbe7cZro2Dsf1NqeMRc1chLuHz9nVgTsWd2FeFNORyJu4apwr
SB7iUIYW/YFSrd2Vdg3c1r+81JDCdB+BVHcrDTozlfAevc1WFXt3PN/Tqv3n5XSS
V7CwwjrmHA4kEP1saNnoCr36JVYEcnWpQj7P755YIe+J1lzIiFPlI72Cpyp0yzJb
dYwA4IHm2/3bQOMAlhIt7nwlixrUp1TZnEZs+d3RK7ITdiWp/97UxoBLSnyMBWHJ
S+G+wuMzkncuNDljPZjQV9JCVspAnB3xN1e1EeEMkYxK+t7pUvdqztqsDb61HEUq
kXZ9c8Nm2uXby6zZg7yr2+kmkQHYO/KnhX2hZTvH+tKLZPOWuJzGq1CA6k77T6F+
FgpZPB/QLfm8iVbZ7LEDz03pJWR/Mvmiik5ltdqE8uXiKKd02su1DllJmTgv3f2h
b8cwSWgDxVYQWWd1OL1/CUfcK/0VNx0SsI1TVfACHVSLipSQCm3/aXlHOBEasDFy
VdSnHsRMKf8JwBGk2PEA75GheyymMpoTMCYwyZEnA4XdpLscREfFMsSqgcuK4ikP
2K4ZJqfpZ2oDnC6zSwuwyvo6B3R9ijvwU7dHBwk8OaXedTUSm5SGCTCniDbOe+a1
rCC6gMW84/aro3oUev6MHaMiVCzoPx5ipBrKNaRPfaNaXPVQ/JU6ZP0qznznNUkl
/xsQUS3QVzAoCYL6niwFxwRu+m1N24IaF399jFM8KokPO8nelGoluKKV9u88pC8a
Vvuak060jVhdjv0oNBEnzm5E9ItbPVkQfoqL79YQ3GG9fSJTiJn1qrMmXE+R09Z+
3fyKnrjM3+IDGf+98YmuAxQLKPlOEGN1FHUgu/p0onPc0qWjDSmr8FZZykCxue4w
L/V8QEnvkvjc9CyrDBreSECoAZJqfMvxH2cz2KrQbQOatvKIDL3v1zUXHKddJOMS
ND3w97aEk3PaUojPwiKqRBa+/NjS1wH7O7eCgG8hn37RT39toZ6pQ8PlNyg0QUka
l7Ogdc1dQ1cHtDH3eU4C5Vt6dn37mxoPY9QceR9GWnMVR0SHrT7ubGX+5N8YwYAA
w30ksswogaeT3xfKWHSxXlwWTdaFwmLiQUMimvc/SCcheaPUgPpdBWP5mTGgs7Wg
ED2BmdCOKR88Oel+2sOn0R1X8TE62Cbau72/JPQats1yT/330YjXqXaQPVYMaEnC
I6MiFEFFr9MDn9lAjpGkeEfGr54rcPqmqjn9T1uDkwkXloJIQobflKszYeoYEBC1
cWYjxMeFoF0s0Xaj/6ld7EOCrn5xR1AiFTf3qKDLn60H5Y3O7oQYlkMwuzyiEiXG
uoT4taKUKjkT0dIvFa1qlE6RkSFiWeaHB+wDr6ZldiGt7eWPqzsAWX4EAb15COlC
P4xpoCXscySvvKy0sPduy59nRr00iHpe1Oa7fU9pqz9EfOVK7Q5O2LiJyeJ9V7z3
o9kQmsp9Evw/lhFGDAFaeV8LXRGOr24Pgdws/ivmjHBvad6SDrt2sRzvXEzI0MhT
oaKA8kK3SdrcDlCTqnCfQXBKRaC0LE7/B6GTQMUcBZNLRPmuS4QyTxFqeCzmj2Fq
I1kbxTfGMwvyxej3oEk51DVp9XU/fnnaDaaiSRsQ6EEjzCu9SIbjYj/s9EqPbhi+
abgc+2tLr4xFBC5H54d2EWec9B9k7ZwbX7wJ9Dh6f015t69jSkHsNpmkPMzlFUIM
MO3KSuUBxmriPkt6sd9GhHwvOKyGUu6KakNfJ25sNULKghmMlC7fXWxq0bcmtKJH
SKkuAbYQEc75g6NAeQMevhV3t0DDVKaitzTgFeUgQ8P7iRVEuW9oCksigib5QfNv
0KnAIm6sCgeY9W4hhCk1K7stF2Q01AIOoqBt3yrZjJR92GlrFVxuQrs6Tq2RFkt8
yMlJJcIHnC1/peYXpXjj2IrXZ5EYMcvOXFAeAqUu8MxBobYAO2Nnbbd3a2aIgmsL
Tzo/wxurw23CARTmJ4YD2/apsKgJl5KfUQe3Er59QGSLBUQj8FrelVCFyWKvoxiO
3fFO6UWdmEGEE8yu2D/TptfoUy9lcCWIi61MSC6V/EfmK/VM7vLc8/ibM1/Cqsvw
wqi9fIA6NY6kIFoqjQuJYwUEP4agjDAOXz1eZtjxlwGNZ+FgqfPORNzG6hhkspJf
KqzMqGbMCnD5higlDnRWquZXXuZpv4daI673by460XjbHV6ycXc5xPWfhxTKQYkd
6fpZTQEz5kXOSfP1EOc5cMMsKRqDcPBe2W9m65Posnd0PMJk1UsEUv6XaZ/VR7Vb
lVf1tdqi+Q++6et3qr86fkF/uDKMZbcmmSrC4+OY6zoALfLj2r+YpolkbJ0LDEcq
cmxRrmsUZebXGJhYFi/6PnwvBDv4g4RkMTSz9eU6bfKjZxd5BIqHffkoO6rdF+19
06/ChTFG3zqvu/a9U7IZDg1sxTsLiMWLrz1HrE5p6zYMmQNakzIG/nCm7swAqZ3H
Js0i+UvXogzQh0ABaNjLuU4lnSt7HgOSIteOBXn60fgukEq346vnenarvBXFZK9I
0B5/xXo3tjtOIVEn7tHDzZ3UGdFSv34FDZUDlfqLtUhv/IBkHcWQUX/34zzOyLg/
maAATyyeWV0o8P6ozdgkQ61dNm9djZIHEwWp6Au2CQbJfElFUXeTtYIUhiDENqiY
RWlzfcZMxZ8wuXQsAYQyMMnaRQAEzUTI2SEFshzeB3KUiSvSUlF6K6M61Y/VbXiB
1nevVNo+HlX4eC5573pXg73Cs8l6mp070+Geuib2OqYGkkjOLiUUB/vyMAEONHwq
AqUkcR+UNHSADjwhmztl9H355uRUpCq0XVtQH8zDfass+6Xnkn/uXXAoFv6jZ2UD
wrT8/U2W3UGmWmC7hXsw68mNEb3uVHlMR4fCWq2qmfCqtE20TeodWA7fSmkvRA1L
y00mUmXPbH/u3PzHW8HFse/tdfJWCcCHMkrF1uuJM3PEjcingH7g5cmKCT1XgG+8
45FTgsSLHZk7GGf3vylGzBsZXtPkX/T2H6/Je4tBHu95N5yronV7VxDUm2pUMtwd
wAW5ucVsJCvs79T4B9Mhl/XU1BHgrKzrkRnCLX0IFjqf1wgupGw5g45nT/DJxkY6
9uRc0J3pySNyM3HBXUpccc8M5eIogHWVLg0H3AFG2sARvnNNVWI2Y9A4QV2ZljKw
/Tiearh1v0hFMaeEJV6NdumhDmkR8LR4G0kW3u8aw0yY+mzqrowwB0vOpw6Cb68z
r517SS6Eqt7wNnqorQrCr9dfbn13HNsdyR3MBDILd87x5aENh3M2eCJoKNb+t+0M
54XKeyeAke9FY0+CdbPuBX3JusOLYGtUgMP/uw26co4e7EH3RpVAQfzGVdKvcHig
BTidElI5qT2Ob5sKtxuDcNOvHfOds09RAq969Yqxo4/k1soy8ZKE04Q379GsXPTk
bnJ1e2LEGw00UUCVb+xssLZHEkIta3pr9eSlaYoDIFS74R+ZjbRu9a04k2tHS8JZ
sA/9ZZOGOTqJyUep8SRKM2h1Cw4X3GExBkgaZG8zFZB0nvHlgtY0da6jcXZyXA0v
JXlGjwpzwOLkXqC7gG6FaOjx6N1mYGPuVT4mktFzF1/+jISDM9TdrjUmqWg6PgCu
2ptMQsdONuF8lgJgVDA7OtDNio32oKd59x95M+JIRjugyxPuz/LqH2U05fsS92Iz
pGHw6DGIu6ZriuGWxiojZ/JbV3ZfRT1OQ003oImUDUkacxL0q0Oiezmq403QiBOg
/eUcMEg2zibYCmpGLOz8oMEx+RN2MDb+ryH9rLmEBdbVyDS8U2mtZ6kwpaoDBW+B
rMyEDjd6R5K84kcaPeFLbuYvGgUOTThMAzaoGvc7XGaA/6nnWr0FipdpLmz9i5aZ
0mDQDRLgWJLvknJnhqxJngwPKQ9L+JkdDN8vAzAZua8675lfJU6hSN6204pS5hsu
vCG4Jnzk4nB22xy+MXRp1Kwpq2lzSwC4mc+zMM8AX99Ed0n9RuXYNlkwm+7+bj/W
L4XqcJerXjMDsI9a8/Ho5T0tGjaXn1Bb4yDGwcUeXmO2XQl1wCX8drweTt10/EYI
0ioI3yKaOBudqq8qChL6HpSsxIC9sd7pgls6Vmx28ft/rzzzn8+XZ/Bi3AzQrSO5
HYl8NPdA7aatpkixK+TNtMPnMVkPT/3zbQ2RiA7A3StFAuCELmjZollYzKczqkP/
vJ9STFDqObRD4yrtsL78kjfRKE4PEYgWQjsecYWMnuHgKNuf/6FHSrB91o6P3ez2
oBhT9rKpKEIKHONjYtGQQDrkWwcSDw3zXzEb8UxHjmorfhdfcAahZb08qTVuuBOj
Ohs/Cca+ITdglhFAwLu6STq/PAdtCs0BcCX0uL9vrS0HtIhS5qVVrqTQBb7YBM2t
/7YuPIGT7K+ttSo8OfzMj4Kov6//g8+37xLwHiKLxaFE1epHbA+6DObtmqkY34Gf
z5KwQPo9EroqCmE3u2R79lDDHYXEXZVDfoH9xt/JxTdqsVcx3eXa1nmFuRJtHCn/
v8OzIA66rRc6OLt2AiEPu+AlMgZ5bmyE9X3ztKKf5M4iAkTPFsNeisvYlLPhYT30
zvgUZbkl/eGoaM+OyvlzXI6e3JmVUGhvaQzyVc/VnfjIGFcipY3k0v9md3qj5180
D8dpr3uCef7c00287VoAE10JGFXy3olvqyRBnpczdZKLnWD/Uas57Ihat7aHsNNU
Eu52aUZn3NlVM8z4uzRQ3eGt3JsvaZxrK89X4262OoQxl+WDMSeJxnfsFrwWKsjR
yf0ebmVfjrQBh+Er1glcBRaGLfmdvnfUQfnw73seVnDtVsiDPWCO+RdGosOKjNc2
a5o+86+4CZfLD7VSQr82vPHrwXL7ZEF2PPOw0R1Neww3OLUSka/zDdpO6xnIV35g
GO73fQbFeQRHwl+KqTKd4jQvm8w8icKy678ycoUPp1oYldHhhmXABwOqPWfH9/Dr
UOyXKrVQCzIlEAbey7yeTH/M7TVha+pBiL1Be150cRTN09Ox0UmUFWWxJaxr4t5E
7UtVx20SZ00JLx2i7FNO3dSmCx5R4fQGgIyQLBeKoeBNA/q5vcO31ZTYo/t8Mzzs
++e1W/QyoI1gecUgYshtgKnBVtP9/EVsJo78QbBolcwJXIr3CYtSqghpl0k08KKl
NvZwCckb/lKlz7jrwXbZRN8OG+ew8gVDfpHxpKcVWWk4k+CPz6kWEJrYGe13BKRU
aZYypDN5/LIMz5x+lkRBL/+vtxVU4C/4vT2vhiwxajkdtEYxFTVe0T+xA2NrVLZ8
lbHQXXzdz85njtEFETVZvElkRkq7Y1yvoyuJ6jiIfv9doxdCDYGDJHMd+Y5CqPDb
ny+H3bNlzgKL6Ekd9phdfk7GBm8fNnTwl7bIpa9d7typD/Wf8wIWGAO23z0usqS6
0xOkoyLfj35uGhrZQDJ+0lJWW32xqsGtwRQBS5HNnzEsyCbHe0c4/rglT1aSBJoQ
PXL5JLQFGyZwJOTNGSS11z08Hn46KLuSoHd92m4rdTacBiTWxHTDBk1oG0vQKQuB
BqU3fkc5Ieq4YYmFTLgcWIQBysKF2w5fNOx7dMxKP4EnktykJX+TAmfVMskb5HPo
4LQiGKaGyYp0JtRP4BzdJbXr7CqpSVNZ00pxokrln753UNCWhribC8wHomtrLS33
gaRhkcJcmf1Sn+9wQofOgWazJ96yxyNydFldS1zZ4URXCzDNb6+5+++StPrkr5xY
8XYcXKydKyDRPTy6RQE2CQM+yVbXm6I4ZRDS0aBcUi18FEAQkDPEriGbarT8b8Nh
r8NsX9ASpmLrvRPabRdBGM3XY/Nujyv9d8FjldP6f7KFvoThCy1ZiIN1p2pOyN8B
wKtZWN0wx62ACp8QFFLu3OrTkz14fakrYNzGVqOk9erjZJ2xEt7K8+YOlS9QmOO9
tRTZPlCeU023yfRVf1MDzVfsN+Pkqhc4+XWnSM4tvf6UI2nMu/08AJz0tWwAHJvf
JWfvhMYEftczaBBkOIs1GG/QNLgRFSSGg/O171hB7h1CMk197lz6OHOCjJtxilh1
1VzRxE2I3f7A8G6RXMiec1JV8ijIOqftYhwEV412v00weymFZRhyeA+ur1ZhcTMf
2qnyMnqucIWQ8UAG3hpWmlojOqrmq6e6KY+RPTtbalKQrGTVYIc2eaMs5xPCfVJ2
TQ0gaJXHOPuw0WlBXpA+TZKlBcV1OekQSyhc0+16+3k1AACMB4psn8LmpX7m9jwp
caPvgUwHqj+/FMa1hYyY3Vdz39wYA1j5d07PkxBCCHHZKawLbXK7Hitg8B7rHmrC
xrUDAaAiDVrteRy++SXwmkO4e39PKyRNqXhoDtSfWd+RFoW8HviyuzlattvNsdtQ
KY5PwKggyXRzeA6b4y6F7aw2gYsKVM5S8wNjG83yojbG2cJij3+C7o2uXQ6TQlly
PuH41U7F+Tjul9WCK/f3Yr4oLCSjtewipb1KMs7/rupBXpzidAilzh/QQGcOq8lK
WWbdh17C4Bjqg9OAcLBttfo4Xme9ffsVbeQMKGjzvtQnXRussrlb1fDgpLAL91br
+bKPsDjlcl7EpLqhNanOno4RuCpENgIPUWw5FgU0QE+aT3vURVenmwl8250y2BMp
5jRdf4pzb4MKMJroi8A2SuF5KHTc2DAslBY7sQOR02oiAlr7BhbkjgxfSNWjHLMR
WdFqXoRhlDBvz13XmLZ3LkRQBKfzilshXvGeXjDZ6XrfMM5DPgrZnGP5JqP8VM2M
8ucHq3Hg2wEJ+MwU4NaewKdLIQ/+6d74sjg6uQq2iK+cS9guoN4hfk+Su3qE0akG
7nghECpTebCJI47nfh6IqFJqasZFMKck22UIXhprQN8hmVm56ccozgufQH5GxHue
5j9xXesj8Yii/uO7Qr3+QiLxRbUFICX8DH3whYCuzDzYHRo3TYkHEW8tdEuRXZ5+
EjM0aeeKEEm1GBA8yWGnWjKIJzthI36KZxJXS+Y710T5WJ1I8gRbLRtup5XgvQGU
InApKQTf5svZ1/xFPpBIlo+p2lJqEVPpX1mbKI0ArCGbPlUm9YBTnhthfj3ebHrX
Gu2ysPPeEMApovU0waWs0qIZ2fkvd8QQFsBVawWx+ZvhNesMu3ykW37ppWd3ZlXm
EY/bqSXb+qr1z1jYfnL3X+qvfqToddKG7w8qNcBnTCyAknTTll534uhP37CdwPn7
a5JH1BhIUmUYxeStX/szvOHxpc2X/cjOrEwuHCfxjYzTRMo4xgZSk0idj5dv9AYQ
fRKEe2olBEEEFs2rrpLXb5CQI+c48/vCzobghrneN8d3ltNxGuNC0zDN8TsBLaeN
cF/gQMS96KOwB2v5svQiBOmaf9b9vZvhtY8GdK+W0f9iaMimYptnrU3b38BVJgt6
+9tHBIpd5zlnQufxmjbVpTJ7HeSUqMoufKl0XeilUlpe5wwHQ6padYVw09KldliH
kXqAVuW/PJy0z+WlXQmnqxkSpiy7WjZg/l2jcCf8du2kt51cOo0w2afe6EriEoV7
rcr4Ve97WUzVopAwMxrnrRUIEHr9OHHCDKadg+9DOVJcj4OGqyVyKEW7w5W4NzSa
QHFleopVCRVD3xqxH4OKibbibZFiFidKFw+bMF6+Z9I82xiar2AYm8+S2kU9LR5Y
Sp+IoHy7QgnI0Xc5LNr8tQFPmlW8aNjXrsDdTDFv9ZCXOXDynjmLaEuZoyrmeSDd
hK+6Ju3ZYVyrFwoP1UvbBWNrnVg/r59qHMuXOIW0+wYL/m8dZGwRqiavrR+VFlhw
dLq0ViTRLOZ73T+zHoAk3BAMklasoCjI2XT4vMn+7wJZuxt4TQSGXos+lO33Yxhq
KVgGDvF66GT+NSOIOkMrIl0V8zPCzH8zNtxzNNRn4Qb6QFPrOOWnCmT9LeiZdIzU
FFiiiCgDkg/dJPHgBcra0TiqWkdC/2CYxkRXntsOll7SGrcJKK7Wo07i1ACwIEpR
xgJ/S0j9pxCPWgxz1EIOLqCVX3Oj+3XQHk9jMZOCSG8Gihi3KUihhNi/VayfReMW
saKe3g/XBcK0N90gbDttphVPYAfItCo5uKTMGYFmlyuTOp5C8/0POqLnnTQClBxF
a8LPApUr/fNuan1zGXYOhzn+qcET2x4Dwn3w6llYE5PH7+dRGwbpah/RxqOD7+99
TNncK5RUJFrO4a+62OSNOULuEBJK62+zYcRTOjf3T6tG/55c6/N5+aKDOSexaJ01
KH4EG/g4Abrq1EcroC16vZhdYg6frZUM/v7rWLZjudGmF7/V5AQ1txbviXfnlc87
4basJP3qW3OR9BvEmxwvSllC9QvMYemwYzJOiwe5gFJG8YWsy6biQbLEBMZaeByr
YRK3FJEeqFAgKntRpA7Lz3M1mX6OTn7DnL3x/S8VYrOU/CP/B8+ejrCqoE/LucBd
4M7BT/+BYLtfiPYntdt9mAACCvhspg+qL1F61HB7K9enhjcN4mQ9VRrWk67BUs0U
aoulZCE+g+HtzLU4yRZK3cEVa2LBoHZNc6wapWtFaWAEgEYB/breSc8kCwgS+3qW
9/slRaFLnu/0DoNDGnseYHBdWt7LpqCdfr7kL/BiaDw67Bkw0j5ltxg5ZbuEh9gB
wcsLnLshw26dDpW48Lr50N94Rji51XD8Fvpya7ckBI6n8cLr7d4pEul5UE/d7A3r
1ms9RtDPtKtnRQPoK3fiDwV4A+548vqo+3+u8H+bEut1Pqu1EzoshsWIVth3WGFh
NRllV2UG2HOzIsS+K9edt7dayXKtpyV3y7GvuRt+S23c91xqGhxwNugREI/IN88M
z5CX7snSuMu7P43Dyo+6q3rabSgrNGzVFCSZeGSECAQb3MxH8AVGMuRL6iBksMJo
hZaeEF/uBiNZfNpWqX0CLR5L54xXxVk3czG6BWDDGJlVNcHHrT8vQFKpSfUU2fs7
jlOfBu8QtgIAEUaLqk0+hZYL+OPBYsX7KidigSy7kOqEwPw24FOBTxP7N7sOiCCt
afVA+u1hABcvFnlISpTM/0b0ggBOluQU3iquLXtGqqkIYr6Nhtl/kC6NsbbhYpF9
14W0e3ChjOub5yMEQk/AEbEpyt/URyi1IiGuEzWWeFbp0g6T6N+mKOKwatV10MWL
3SNO6KvajGc6BwCAx7HqMM748m6jJ383lJUGG08JKRfn/ND/q8GkpOwDNUTJDWRh
KvUQWxgMAkOi1yX9q8pNcIkIXeCTSi6HUyk4oQqRJYqa5VwLl8nFzvV//V2iilE2
wFPkCj8s2V3LBcr0xXSzOABvBAZb5hFamQ+HnrCUpH1tO9yxh4RDS0/xddx1oTQ6
s8aZSM24GESxGJ1xSF6QLphVe8KPYXBSOhsspw9ymnYkE4pKTe4ZVvsHPD59iMHq
Vm5kJxdg6+dp5dYabCchBzpkdkFijiRZ5dOJPjot6dSzszi/sPL1hXOSaqpJiJDh
YIF3TMjoeiRKqJv7xMG8DifVceDkfFIRfdXOQt7tmuYOKUFY5alHJI6e3PeTFzlS
/dC6enruBzbrDU8L80qVnjw0Dioao/ZV/6WeiKlB/3+maEhr3RbLfzm5Vup/Xgny
BFvlO9BDsOEIQXkFcki3reBZgGpSLPSnKr/AFBAbnTY5PMw3blmt8NFhMAAhjrHa
8OqCkgYjfYxVEYDbhYamdFZ3fda9M9luaSAZ5YT5foJcyIiIJmGwLiyS09a9IFO7
clJevJWKLK4JkckIKVPQYLFq+AOkXKoFZ2HqOxVW3Q1w4ZDacNV1ZPjN51rNmDBQ
/rJOQvFEwkScOlPdwG9KF+l9xhYi2mxAevGJRfYRZeUa/ydBrmV4MMEaK/oKRC0v
qDP2zzjsSzmMWr8pHHtMNvIFGsowcKnbehWQ2XzgS8mSSOvoODoUAooAvkqZ8WvF
jSJFn7Fm3xxVQLThAGI4e0ElmbP1xVwo9WUjeE7Q4wi/66wPGU75kd7Ey752NA2x
EDCPB7tnyqraxKXXgVgwTp8s0rxbKiQ7movNshlugA0Jc1/0CB4Rlb89wPg7if7b
SOZmgAPkSVy1LXqSony7am3eIGz80V6/e21Vz55S0nxepXCX9pA6SxWuo/QB70Gm
0pkbcZhxblYard73MSVIss6pohMnLPwo5mTKv8oojM0Lr29PkKq+Ygvvq/dXdyoP
G56RfCbRZKxhq7WVcCJgDKtNvPKI+YDvzrzJ2PljHmQQ6ip8MO8AvQPm0Nidpq3W
WHWS3ffHnUb2KirvtWZDSe2KElO1C5Whds1UFakIQydx0oGDTVtjFHBkWguC74Uy
5kpHDSATz0hvyOVHmemRcirBYO3Gef19szaV5lBiUdNkvpxrQZsU1OssqulP3l5b
rRnqgwyDLlD15cbUiIAC5Q/r5vYs/2JjPfeY6rVWkffR4hIS/ozacCzAWdEcrSdi
w7KPRvvIUxCClYc5C+cIHzsAcm7wdz/Er96Jon7V30RymD6dEv/P2XReenX0FdAV
g82HfaftSyQh9nykLRkDRwVs5hg7JgjX9jUPvofzBRsFqPOzfODbXXvJsg9mAr8q
f6Cc8NpsqoFXk/pUzNns/eQXCwOZ3rp6w0fSUocp4BaDnZ9N15D79G3OeAhbKGrJ
u4FVlPx5I6sThM/LZGa9jNsk+rrZLE6WoGpeD82z5LO9VNarqj5YdsNxRgoHY7IY
AqG+ekdtT4wTWaW/Zh/on8vqCaYA6WmU0wl4SPCOMSz4xryPbdvnFfDeyT8CDFWC
0C1vd9Sp/+L1Iu3OMRimQy7/04eR4B23EOtYATtpCpsNIexxEGmKK1nKPpJR3z1T
TlVD/3m7wkVUOjCkwS/fSxddsbi+LaagbtUfLLGUvvbB83u5dM7Xtb7JmEgUfCN5
rnKP1qZLoX3RAGzQ3Cz3+j6T/DeB0qf3D/w2f9Fmp9/S1OhRPlg7GccgMn1fbB0i
E3EwdQetODfl6H64rivw1KyHoJx+Pu2er2C51w/VhHuMLA8F5jUuY+VIvFMtPwdC
CvsccOEoYgb625AmwKy1819/hVFCFnsZuWeRCYO0g8DvWr2fpNYzum5OnMQRTC3E
YiBzE3afnmm3D5Bd34v19gIF8k0onAqRY+E1khOoFYOtZu2MuNryZcvfkHbtDv70
2b1rFILBJFA+zpI1erqqkrCGM3Dje7/W3p39m9tE7e9jxPtM1kgOSDa6E1S8RXCO
iTq4ptEOsTIO1wHweQG+UZetYj8K8/YbZ9KI6iw5V2ll2FIM86coCZsQ1nYHIIa3
aTVldE5jLLedR31mheCgMN7XV9m6OuBLi1WYVgsZKtDhbJwzoO9bVTqcG9igCWpN
tvASWHtfK9ZPY5T0cD7lM5rwOV56HTg2eDlial8AOJNeLD2IpUQ4lPsPsGvdvKpY
aypX8lqt8TEg51LQ8FVsZNd1Idx94W5VPjfW1I/kuv+Six+OUsKtGvtIVC0ZrFn2
lhEZc3EbbseJ0kEylFYB+RkW4dPVhG2dqXKi2Rn3vS0zQLAfK8rLsgRSrI2L6kqD
hPbx0UswUQvm2xgT3iPgCuVOFglxrx/ER6/11JNWhkjPeWEb5wjCK+3P1b4v1YMw
VocKWr17pxJ+IDISR3ZT/rRlbizChBdCD9L82RYM8ti+meW2ZhbYdsVPkrZEW2JG
S9TKPQmS5HWIdRkHyMoPCs0Yp8KCmdNFeZByvQ20yyH+GzMUNoGGTOQ6RRwY4bCL
mFUyJ7E4WFu79EXrWnnDfhGG+usk2uuW+IG+01Sp1oHZyQAsBU+oZ4fAeEHsTZ6l
LL4s6+iagsVBCPDMMd3GN/VnFTdeuZy6EdbrKW5ePtV49Srd2B9jZRgM/F4srGha
CbCUAFt3fBhpTN32l19neKE3srPO0KaBvYxb90aRqI5poR8GZyeGCqfpjz2ECb4a
BexQfrbFxYSlcLx//Q8ECJrmGb8/kd5fjrhXwBPzp79I015tajhqanJqNDDUW/CQ
IwGb+V94Xi2JbkTXWa19dI41tJofWoXutjbmT2YpQ0+TdbWQLeORlMSutRLQPmoL
imndV7wpogeICoB7uP7wNS2k2k1cLcEyOCL8gyMf/CATepuSdQeKphLjDg6ag0Sx
R0CZZufcA/Mcgy0NO9AXs67vmWnJFyaytEAUi07cm0fKuW52OmBSkE8HM6C7P3HE
/leT4sSuk5o7MFzjonXJk2nN8iHwFLl7NNxvYmxH0xo+/C1F7PVD1bIeturdUrxp
xYD/bnQuf4Om3PLQae31ctQyCjs2ZyuhaVq9UWZXaskgKLRjy5uz+NP7r1kroR/D
6T46Ny2gsTWy/FJGmuRgDbryVSwmI0e9odBWdrA844JUuilFOTrV+hrDkuMNu13I
pPhOWALyQ1I2m/t/lP8ABq+GD+88aZ7LrpvA88zrArw3d/TaSrf/REZdNeDA9K50
CVNIKYdzUqizHnGubuzU0wGzk7YjgtfvXVsUkdKqWirlkHCXbR8D4/GqgVDr+IA7
KvfCKvoM6+UYMlzYFZ1btA9lJLjwEXuh/7qhzL3ZeCydcUfco+O1p4iKBUMnSyc0
LBE9gzwMLD+nh88IAjBYQq+PJAwrZtEzxJuuZ4cSx//Tw11pL9EWqodWcb2S4a30
h/++Xhge/JdrCmCgygCYXQMMWJvieQ5Mhvz+6ChzsacKDpPZ77/HLPSQ77zs2bmt
nFGofw6JAGfiY4XIJ6lopdEofHW/doG9cUayJRPgaPydHA4ot7TVTY0L7YAOr89b
1in1/il5nrKHTF/HX7LByGD9dVM2eiDJTwfmkBeUkJBPz3im7gezWqGLOP2gmqC6
6zVprjPM1vQhl8tsgU8LZLVzrE2MiBtgu/gP+PKEMP43Frg/BpqBdHQNTBco0m/3
qvDIh1OM8rXr8NFWKyBuRgPnUjkphSUz68ZVoEyfhChWf6CioOK4FV/23wO7z4ku
hWIwvCUxy1P4LFM1ReqMH23HeI1wSmts1Ne26XnvwrUw0qpSNco0nShlYAh+uqR+
SAEuHac1W0lbQnYV3AjdbbdKrZ3dZZfUGyXVQHOvtTAzcHBfFQwPRrD3sRHgOalO
u3CKeJM9Yz14/wPuovwLrCF7Z1w9XLyco5X1d/L+IZ8HIrH6wqw7QZYqNRbS5Ipf
4oGTlp8EOV80rHghZfynltIpofrtVyCZb/mGQPJ9fTOOksScHqjnzqVvD3dl1jb3
h/w7zXD4G1EyIk04d/qq45ecR85/XlenVjfDCJw7gGoAVsnpzUZMIpeN4rhpbDjQ
bdTr0JUKuEtmDffUSQCaSyCxEGH2F9uxv/t1Oj9DuFXCPL5Cqlttg3nYw4mZotLt
Shp+c57zXiCKzJOk1YzoBeTc8E+Z/FZBATiwpR9Tfh2d5+CG7NOhf3wJijolsAyY
g8aj/TMsbF3f9PpuNiyRGspG2y9rY3FyqWICM73au/MtcsorlQ2+3NWGPTJD30MW
TmPrDvuZOEFwJ2OMTfUlOzt/zwHbhx/gw/obSffUuzYeyyd5SY82cgkc1XnMhPat
r7DmbJFScTDts9gHGWgQpGKN00f7VL0Oei3kmNMqLEEsmEJcNUGRdUwnTkK+z99m
6qwd9f7zY/C2fO2hKBxpuSImYgEqEy2dz6qne74eBw922dOwVfa5XoZ3ofecEuLB
mGonxgR2fmJ6vxb/8IwaGKPdQbgK7HPpfER8wMXLyV6M+BQt828lWaAKPPgocx+/
aEaun5k/xJIcxZ1+W9REdS6ZCcumrsDwrq17o+YFVjyY5g4PwAygcx2Zc8SwW/Uj
MPmHYBYcXm0OaerDY5rNNBfSocV+UaiN55OYAGRWde4PCl3eSOLjIb4tOgHGR54y
BGflsQDW5xQabarzeZdbUR1CGXm14IkgMZ1I/8/Wyioqolmcq9Q2PHXvaGOGk9ap
Dl5u2Nrg4na+JUqdY8rFrhQ96wZRnU7cMlPLiLaQZMU6RXOLSPNRibWyXCA6E+nz
Olwq2FASx8qv3qv6LnzIKD19aIz2dqzPIyKfUkcfx00vZK4HPoQ3Z2QWjw/67kdN
P6gf83D54LBO/Eoa5uLwC0KRzbDKHXYnUP3Jkr2JXY78icaLbKEZYDYUrlS61zDj
2R2afVHo0uI1lTve4PJ7rxZpbu8y9yDPfv/Xb92ao93mwexXmgtl5gy07P2UN077
55ktc8wLqKvYdFmV8g/18GlefnGn75FEq38xjgX1wrAAO33bvBY81fmuw8KFouVi
EKsvNN+gUoMXJc1P/J0Sk/6vTYTXl4fTNOtkNSrkz29gAM5JtAk3n9RGPwchYBMi
D+074YmHQ7iJXcSINhzladDslI4ycB7afdwupHUpYLY4vAfrD8AsDQ/Dug/piliY
U35745gFw+7I4zlyZMBAQgPXwV1UnxEw1ekkBV/b7vgL3bnXKmQrNp+rQLKdUq+r
DY5ypxJfq5rlLTBwfkS5bNB6/hmHZ66uBjYEhELekkA8aS+CY1GQ9Ypa06FRh+Rt
7IZD1ZkPrKN6u2JwBfvYD5JfjD5erMzMfWpRWxY09m+JCAoLJb5F6YVQJ4B6aURH
3xsfA/a93aaG0eErqcSUeMVEP4xNQeAQB4qdjMp3cacrkm0ITfjyCHeyMCYpKp2Q
zwEa3Ni79QS1o2gAN+YVpigbV4aeB0dJ/DGjzY7xx64CZFID8UStecu4OFBGu1Qn
rMCfXH0mvcvpHqGJTzbnRHpE5CEmKkEYD+uOBCaKR0SI2N0KO4/maBigfgIKprmg
uE9f7PScJpBTi5H9m2Wn5ueeNorG8VMXI6kmeJ/pTzNW21vdFyHoFgdinfSiq7gf
QGm+rr0DRCGXDehI4bdzbMM0V+clWVESVqQu8nuE+j78ZBGlsREdG4UrPAdHpmuR
fX0sFAgV9xL1fIGeVF+XbqT+cangKEx5al6tYSEajvi3tZ1xi0OrmvowA/+BNT23
Xj9n1sRGDOPkXdai2OG/FqZOBx3ryu24D2ziDqY5nJ/6igmpyYPeB9gwKpbYRphB
eqS3OK7m5K90USQgCWYuPqXZoq8HojDGHKoz1qMz2UyjxTIpojR1fod2KNbmNFuU
Thf0CzhggYIyOFI+8pmYaQ34Ll3XAGDqPm/SbXvwHlsWxUTRE3AktvvJm6APieOR
CHObWyPqxC+MkbesiDtKutccFZM9QPnjxD5SPoynds6f3UK1CSO/eO/Yqkgdxd1M
ABUEoJPUq43Ra2fOyvD0RZitcMAZySXIzM3IFyKllQSZShdGyV03y/TE/WE/X7Eo
Xlae5FMZ5Q0u2FjCp9PrxbUkt7CpmhzevHW/u3K7bnnF44Ne+fWqO6usXXHmUGKm
oxlgElb3cUdyT2FqljtZ9IPuxbAZilTb7BgybNQo9trMwsOHhQmj6Yk7t851yXWr
fH1EIDct9kbcKIW9j6ESpQ6MMTqWvk1xRvPSvWoZNuG5uX/qCA6jyjlCqyop8W1B
Nmig8sOIxmYm7VYxYVRBpJH/q/Dj9WZrgvhJYax/xMXKpMypGwiSZt2oBOCnWXPy
2AWJiXzhSr8pR92VZUxlDxTBZCuGh7ODF7MOyyrrsQnHM11N4fMje72YXbpmoxwI
wvRZXqhaeTtBhH5cM/AjreEjPxCjxTmXh7B//CDPuX/PeWiSyz3JVnyMCIzlZC+l
6eqnuoRuxrAcC9HOLJpVLdlMlgjGOaUh1D6hy2lhlHAQSPamTyhlmbv2KwvAvatB
MAU3A5vdR7tjS23miKnrkc+VpF7xEZRXCodsyds0ZLeV19LZOB8XJMZ4enwGFjW0
QqHUSjyHbZtzp02TJj+4jO51iljB1SlKPMtzYK+vZ1/87fE/fi7M8ojUEtNd5FgT
sFx4/9k6KR8sblszAF6vy5InlZilABWRiVFHFgQBv72lplE7/OXB4/iuPYndXYBZ
II97XntLiYGou/owq6AcJDSoGBdFt/I7wcAAosIlYwT46TwIPP9sKu3YOaSUEb4t
Oz0qizMhDDnUKHFDWjnSJCIH+nDmTqGk4I1FZfBLabsnfieTE/4LxodadJmcWvN5
UvXgizg0tv4r2oJ/7l66yZ7d+nYYjCO9udawG3azyIF1KSgtqEQFfQT6Z8xjY6A5
B3TROh0TYfK75ytMivzHjEVmHcW5Poi+pB/bstBxsiKq5c5f19PV4ZPFk86TBLP6
nJMsFQ86MyBjPA4GKXMRDlfPRTKop/GJhdlaqt87/fLnkh+rFqHctNmsnos8b7mC
xwfj1Jm8bIBFXZ2w9zcQw2rde9rpdqXjQb7Vnw3a1oOPQKZQyq+syQpem9kogHSE
KstEwbyPX5v9Br/hRKopJWmLVL53/eS92lQK7jXNo+KItDxV/0bPfsUVcEUEZePw
xRgk2t8LnE9Lo2rfpKMFXmJbsj7xOiOBnblZGGNbGgYdRa4F1GvOMV2B40pHGKuU
73m5xze/U8tm2jnX3AzsfXb6SpNMjDvsG1Nxax/aeu3IQlVMBCV1V6gCs1Sf088n
B1gqd4czIUHEYHo6GiuCYkVYnSSwmkZO3Yao+bviQbwdsyQ4ho9kQeMh0gQCXHjL
+ew73z25B2vxEal8iub6v7XKBlKnHuhYDR1dLgZmbyUlh6l68BNxd5tgCzWSGlZD
yl7VW7VI5s4wF3wPqFBXhzgXsuXcEnDBjmOEcDbcQtQ8lln0uAo+yX7byAAeY4Si
yhomgbaUOXzvBsf2+QrQ3N72WRlE6G1Ex3V9AS2NWwd5E0S7v7eQCYZKgg6COZxO
rmVYt0BDh4iGMkc4TMxwKyyOYKkaKj4W9Ju2iYe1MApNCCi8q8+is8qRdrpZSUGe
zLkyrWP/sfRDJZB12jOSCtnZXWHAZ2c932RC3FRT9ATp232c7/KxpubyTy0Bz/kc
bKvnW1JDIumasUH9rQwW+xi1ID651eaM0uM/ldpi+blT4T9rCd+DWTR+Nr1GNz0h
7/soAGRQefiEALkQyugvETFePpHOQuEPFBqg7A85Xi625DfEUFqYfEcA5DyyqSZN
TQolSYoel/W8RqIkHJp9Wzwdz7oxkx1qBK9dLlTUphqVTlJ7uXDeKeKtv91y+Io6
QNX7ay+QYJ7LCVn/y2jtsgZApTe8rfwgdbY74hflCAm1PD7DPiWxwl4IfyeQa3qv
CHd0Oh36cusKrWdEwSo0k9Hn9oc9qzmObMDvIbxPfM2zBuM5V30iE2LjSvKSi6Np
tbS1RlrypsEMm+qAVmS9G6Y1G7hB96Tq5qAVQIm66hqS4/h9yPczd+6Gq9/j0CJI
bT+d3ZlMSMfKDgn5NdRd19SgP3+hPjfdCzchF1a45z+KGom6FKzPjDCkAhGYAOHn
HbG2/ewuXrVbdIJSSQdxujtv1FpVvn3qlin8R91uXgpLUHXlfxulkOsMmTPLBX8V
JhPXKBhD5uirdh2p++sOJfs3wlVirQFN4OgKgDck7hAaGud4nwZJZAtyG5u5IXDM
76lKLaB0UrbrMpQgbAd+sTXM2mGpeomeY7SUBk4cMWAhg9vEO3JtjmARWaSaOygO
zdx0CD70QsWdHLdZoMCtwsJjk2h2ghKlDQpM3ekkShIdC7f+MdHetFCiBoBUwtjt
V8pOkp7QLdjcPtMtT8aTGOWTCt4YwDZ5tzn+zoqHdyNyb0ang7jOdinI38Rw+6bT
vSprvl5E6wYNnsvqEcgbiqZS+opNJCfukbkwTVJqmng9n/zUcAalIOveMtfx0Me2
DF6hqLcaNc71GmUo5gugmVxe7vLwDUDtvkSJvZRV/JKB779MBDTwRDW6/54t1zMT
wiUvbbM92rJTQ9ki7aFc6p6PuhyMdWk9nbtpU0LJ+GFJiIYVtYB2k+mYEoVna8Ki
CedHN23Q/kDmlFavtdrIjW/ZlqZNvt14PfDVz0V9ZatodJo543e6zmlvRalUqZdW
O4lxnfRGtzm0FUlGMjfJL3ATGYwCdBmDL9piIDIW1L9UfbCY1FI5Zakc5DBznYlU
nR6fIuWU5ctxJki9FbxCRKwdo0JlHDl8Y+u+1oLbNyz5IoZOZK+zKUQ7t71iJeuj
+1VixpjUOHuL7X8RDNQSYApjt5SEj1y2dq+UzoaVpFx1NMfeZrhQ87bzLL/tafC5
kUPYMD7Ivi57ezL4YSJcFl48AfqIVMHt6oYOgnuTq2/IWxrhOqwxXumeR7Q8ZwnV
HIUjYThL1JE8Ii4Vq/bRSOPJX7ClO9pGqymnXVJAS1bw1Sa3dLfIArLRmzk8+K6Y
gMEJf/g2M/jHrqGNT/F2YN5d/pONw5jiwMyrl/hsklWMwOme4g774CjkxHjlNnfq
aFcyqTds7CTdLVr47cPzU7SijnaQP9gBpHRNrISgg81GN8j36mk6zdPMmz7547r4
Rcftn+Uftubsz/5nnhZXC7J9+lXK9b96/QLLCm2OUJ88wSX2unIlvNH5cx7oNCKr
h0FhaIjWCUxa26pclb27wyFvRc/KssxTqHyJzvpfLtaAyo8MpUiTgHzqMQ9bRYX2
1CLoD0J0nEEEII5Z1OvbqdnAP1rJYFvEUJ4TLs+ELmakUXjOKI21aGWon8OXSQiQ
bjhrBtVz+hp8PRtckhQKF0CJSPJZDqwNo8T8qJw66OC31Wrjrob0JPLruejERAGK
g3PIqg2xapC9oOmIklMYKOGRtHPvquqh8+JPRTrY38Nr+hFBPCFxbw+B6bSts7xX
3Y4bhTr/hA8y7g3jMhWwtBr6i5NmSKH7iOC2Rm7EdJZtqUz/uvQcZK+JIYlK1OaS
ahoXDVxABzj3tTDI+8L6IOABhm7VwrlvwQv9UoKsM0GIvthteeLhce32HrsnpIZY
2Cqv5TUY+3+6a99HWujoAVWto6C0DZXmHDmJXE4AcCPIKN4sh9kuFZPtTYZ7ZPRK
m9iktNvbkx0pE6Q1tKcsAplw70qQcJwa7Ibgog3LQ7STyxUOtg45+X+s14S/+OT0
R1LSFcLoWdKVrif3sLhIiq7lsQHeYSTuYrmzcpxXLftZn6GHAKAMzfZwOjUpjZs1
lqAmbf062XM/GJCELLyMQJniLMTej1OC71vQAw8QMfP1MkpfvqeBCp0BoxZR9D8k
08wx6FhPbBP/SlZIQjnlr7FSCMpxMQnAEFOV3fuTHizXCQ2Q2+ZNlO/Yin+Dr80w
mLR0kafSU4jH/0xuo7ZOuAkFh+tOejK8H0IHaCi8KG8q8QjmzTqRVoNsUKMnRJ7C
O4eBWf+6ErtprWXOJTPcLAkpmOs/sjjUCbolERiSOKfQQ1y+2V7F+UUvYQJFBess
tsDbFZlwuqWR2sFsJSqbHeerfDS2gLcGHcvmkAXRvCdaEmIoqeYJQgI2LjOf5xD7
WGYL3P6aCNy4U+IbtuqVPyX5gE7yyxuLGaU9DIzYbKp3JGIkv2InaRk4QGQfCHtj
MBDwxN9OJd3ej2mwG0sed1tFtlWz6d/NAEWRTBYSFELQ8Cy8ft+4tiv/Yzjx1c+5
iN7cy/rPZZv/tDNsXLsfCJ3ML8IScufv5k3B+m5Vy7DbP/Er/QuYV8r7Zzk9XXSR
RvOIDtjZYOno/fjAJSFytQ58HdVLfmGTxYCqtR4k/OF+J4GGLxHb9Ln583x6uJHl
SDjIZeqAyGgIi6eHASg0OjYYXE3zBpNjMx0BhHFiUtZJzbc3patfRhhSyNUmYtx1
SbkY4jjttbgYYQ7PVnsOEs3KnJ7dACZxTg3qsbn+B9desoF6xTBps7hTa9VWMhn+
cPzjxJOZUYRADK6EglIlccOI1tfMXYZK+Hb02Fa9guNHofm+3DG3SYTqtgZoVBar
/2d2zXBJQpRsu5ZSfzAcmUtH4FjyW+rGJx7Ta2ZKrQ1MdW2ECvPDWgYKpXpbg+3R
/kHrEMmpXLzK06o4nNRKCK4rlRG0WVB21p0x24E5Iy7KmWmJ86SH38GJl1ObKT3Y
9fyAf06Q0uW5W0TCpK3pHrYfG/rXbNiazvQQZZe4Hx9fx4mqy/SOPqoRoU/+qWPo
GRWE9M8vUCcvrbInttz30wS9VGuS25a0rxS8rgKLd90YDoP9WL5D8ITdk68LQhQW
wm8ZKj+oAOj3J+NvBJckN8uLiRJyoTzz9im9DEfiShganTVoYPScJZYVX/53RpZw
Qr30e+GIADjZNjo4VynR/CderyjhNvUO44qLIjLV7RrYhek4oMe93fV19b7z0Kgi
P/SH8MRgDTJZMVk+rgYbQvoZqBGuqRyDRhaQ5sIRUejVwyi4mzpyLxgr53X7Ceia
O5yvqfTYAHd7zx+3Qphxa69d/n5389YeoKdbGjoEa6287UfN6jP0tpJr/OdrgqbZ
FUgV4MU6+cy0zoRw7igBp7KW7GtLn8815R7UvuM18XPGOUaIrnsKzOVdS5WyCY3F
W7psht3ptn22P4Dm5FSdR1gULG6gqNDqCVvBsKY0+F4ZSRk6PLJq/zuXvMf7qCTD
STRuuBFX5ACXxuTtm0GAtNQVpbZCECAUqWCNY8c8OdmZ++iSnBRbdfc1r3+1YT7j
qtVBjSrdGYpS0mqI4gPakrjWCq/mdjQCsbfrxyONUThKv8qjklXObAuu+VpEQ5o6
p8xOh4oCCcQlBONBzN/kcWNZw+CbgTLTu5ioLO54owWhSUa+xNG4JYpUW3cLq6O1
JfRCGW9BrgE+SSkF2+HkfbnHBb7GH02TyY5CWC6LH99vdjswzBtmRMko+x36sijb
XdX60/mNX09XXyqUUD9K+x6Ctg6jJ/o9BcmCaem/6R0zzjv5Ue2e4W9g5zAWwBuB
WEaPJU8WOEYr4bHSovA8Sb2fnn9Ux0LnyMYCZ59JIVfoZYyI4o0Np0R4eqjMTZ+E
qh9t+9rFjyAmBoyJmAKZ7YsjYpbUP8ixmEO9LaSHUrDgpWIFC06E+tcuxM/TC1q8
NYg3RyJ35wIaxWwWMoiHDllg2tqu81+kjRbt1jd7koYPvC4J/3etfhSTSLp/VMV/
3KhiQk9Ao0SPfu9nEEUd5Cz+mzIdyNSZOMtivpq+nYfO8IyrEJ1VAvLierHV9bww
Cuok0btgB+TP9g0MAI7lqKtBlFGbGmi4D3ya08mr3ExNdUvF8B1d9vDKjcOL9OZw
t4OuFFQukGt0DJOxqHll3wZ/Zt4tqEj7tkKmoQNUT+XDJAYZD35sRC5SnG/Zz/Xx
N8FdquSyl0Az6l1j86oe5eP0HuoHM1l+6lwf8PxNluM4hmMSMBYtT1uHdwin46ju
seBCqfff4gVUMgbfZtfIggYb/ei+TL0JYVB3gXcrIkwxju/BNCd6XaoF9vKW1vjc
1v4+LCml4yBXaoWPdbsfUysB13XD1teSMiETWdAT3KaJLimSNou7MUWQEPgbfgzj
EVYRnlkEYD/Th74xcY6ZqlgBSVzbvTQO2MkbXQQPl6JeKS5RxjyoGejQkZuDugYR
l7s/I+Sg9TNZ+eEdlcDe7PTmqrPC+T59yjr0PTnYtGUrt02ex0NRfGYFliSvI3WY
Iy2ulhgZVQIxiXv0h2LAn31DEORuv0cNGLRExmq7V5qB9bCZNNV2M14V60HgNk79
8IzreFPITj1le7VotV28Siq5IcbJupMgI5GRksX10FG1FbA/VWlYYTeV0Ido0aQp
/YSHslumbcJ2fBbTli53Q9ufQA+Nt9lerzoH6d+TFZihYpztb438BrJTI/QXGz7u
17jpWlPT7wx+XrwLoPQLHFg2DiVfzF0LL4dyyO8hp//hTTXnGqkubCdPtGR0M+xH
+G1VKTfmhFhw4Z1FGfYwKxo2vY2lFGZ6vRROWJqFP3pk9eYvkt5HkXk0mmIIm+oK
wdT/Q1aRozYTXw9ImNRbzYJjrtFTI+jqThGRDTWU6uCJal4GfUXTe4CucyWp3HwL
g+xoMg+sEdf4Fx8yK7oFhMLeR5Wwlh57lbl1sDKpiqo7O+eAYmyIzJlnmfT435v3
+zi+dWlDiYP0NWd1PjZPaFbb9uQR4o0Kgol+hsfYTknAcE6hEjRtpMhg1xDBAiW5
oNTYyOuN/btU0auszbhqm7tff0Xz7Zn6eCwpEBmltv07QqgCmSZondLydvgp9fc4
u5bhMB5sMcizb1y5+TkQ/W0CElk9CciSkhQrQj+cMujYMqGXQDS1+oQbwJ3wPfxF
jsg28Rx+lvQ6v9eIB9EP9TVV6MkqVPEAAUMA9E29PLt2YLDOb5sII6XaAI2Kfm6g
NPwujXO53C7LBHAZaSl/Gm5i/kfw5QMjp4BKUc4n25DWctPGsiN0ruBkRRctlAMc
+9JR3RjHM8e5c2CHvAje1Y83eepDj9nUPthf0meNUB5K6VdknDB2jns+aUznENKN
QBcxxj3M537v9oGPfUD7Y5LdaaU92jqz/XBWg24tdqTQBovvvMIIvixVz6+kdo41
evOYQCAF/LWSlABGHJKt2UpG73WC+h08ZX/fOmbjBbugAGx/vbHq4C18afM1SMe+
LZ2GicGvLjuS1DFLaFEsLVPlxFgDpDOQqSwX+o+t0F4lLrZWQQzQDNQQKKStzp8n
GL99qrXvGyugn5nsbZ+LP2ji22kijuwRTRatKj0I9i2RgjiDuDLO1gQBA01nytyS
Lf/aC7l/eODRdU8wXNp3hjmtT+FOV9xPdW0vitYGqwJNlTKCEwtQaYbHcq31kxHx
XnZMwbd+F5XuwUOu+kgjWiYOpnnImg4TBZMiinvxqxlYF3kRzFLXOpECKqbhP4yS
x/DQf1jvdaTOitK4URzIxZreGd4OfOBG7pQVjxgzMVQ7juWN6N45dCXp0IbLjOwH
rmZc/YjEl6FVXUPd4WW0p4qAIEtI9KEr73gyYH6pqRRFW28ddlxR4/NFP4njOrIN
zRUfbkX2iOlSTT743dc4WzoAgSFzb4pkW0APo3lN+vG6mTk51E6lRcKnsGo14rpk
8OwVp9wnpiHVGO5TtuAspPBcs91qw+HG2U2hAaEPTIWy54c28YZFYdSYM/mj0Jkp
cTtv2XG4hVmWFtjP/NCMP47V5ZUTNP5gu41hTC6h1+3Uz+x+MoTE5JJkgLsFgb4Q
kRM+9Wzlgt61UypcWAKl+dk/6cVsCOj1++469n+9lsmfX46ZFkAYh5VXsHm7mU/5
iGxt+ixGzNfMmJx2ru/TrrGjueFladP1TNw1l84J1G7wUTTSEbMHVxCPTgqj9Yn/
ejiVxzRag+kFZOoZhxgCf2rfqomxfM+saOuOuyF34OcbmQXb1v/d0X1tyEk5mHx3
QSYvJRokt9ZcP92CtLeBqj1Kd2P0Awh0d7WB6IiSBhi5mth6shyWf4Bpa1mbSOi9
9TCPFeEs0SLm9h1rk/BKzvA4GuySQe8HiqiA0PmluF361VMy6Xa4t4ax0bPgKUhX
JSf1FOLACuBuO8wXPckMfyRGC+tFQS9OcPRGDSHGtsCkmOVKvV/WoymkTCeLDOWh
IjDM9MaOFoJzwakSQ/p5JQX3Mjus+7fU5jr4P/L+85G4fCctGrZh0pigp+mWvY42
4irToFLpBGJcuhuI6ftgKWZa35P50CY5N0eriHy7UqGiwSmVQn+898y98biaQSSX
0faVai/Z1iqsbFz1vuoZFd8gLyZIZFtN5cc/UG/fFsNuq35R7V1kH/4rhoLK/tax
9G2NZhqNgmmANZmps/rxNGQgQILO4Zdv4VAD4SCO5e3VzNLYIXRHgNUeivwhWxPA
OUUXGZy+SeVTHIeVURKBQ6mM0ZQcXBvYfUkOv95Vj3DTWnKrhdMj8gdK2TK9KoS1
/A0Vz3BVpLR7vUIGAymJbzZp1vArRoiPRsME/XTQE6lNvgxugFVsLMP+9x3LFlVA
C2sGmc9Or1CHZxlb0iNBbg59dCkj8mEo/KWYS3W+9od7mmZ5OgEHm1566Ns6Sf6h
UqLyqyhuJ5tQFet+45E9/jpQq83+hFMWwpUhTx9AkDrnnL5ebIHhnqJpoety+eRL
kp95DidfZxPJVbMvbhyho5c5xxdnW0enOrCOd2nTFvVXwxATP1FMHIEU0NvEQ1Rq
UEVngQyd7A2Jd7OPQoWDGrzB9Vlh8nsGOYw4tfla1YzAZolc6QynWUJskEvGMCjo
4WfXKo4075YB04PWJme0rRcizqMAS8X+VxDvQUIreo2t0UMUB1uT6NLCPIiVczOb
7C/ikYPOxdWLVuzYyjeWLmmMO5CkTsrO62mePKx+F6WyAMcY4FA6ngkZ+X/dPJHc
TxlcQ5mXAM2Iqfm/9PXqK7MybceGd2nfRTfpfecLdEmlm145dB+/eosM54svAuyp
4z20u/Odl7wJCkkDmRcq4Dl7L9r1ZUzxiXX0wQgHM9CeJoyGQR/xc/s7r3TsHDIL
zVcJtccxrVjAiKsXIssZPLS2kljaqApPFxZVHmI0IOn6nMo0C1hB7L7eWPpJ3Pmz
o/qgJXkif+bl6Sp/aJ/oie21jpOee/twpYtcQUN7aY133eARrqklsIBXPHzAjWo4
tFZODGUm6pwd5/I1tHf9eX9ICvix2SM8KGweC3yWtHDEHxq0K1rEP+vTDIkFjo3m
2tkP+b06juzO3uGkZZYOLDisXqqun1vNjYqR+HaTWpxGlyA3UzxsSCduMxHNCbrf
Sd11YI3qOotOToB9quKpzLIdBeImhMKy+B2Lwg7Ou2cCDxywPoWLT3UY1+g7LouT
/lYNa1u9BiB7QLFlJOt7UekxkKo03+LD/RT0fDggYjZsPSTGo1lUB8uzywcxwTws
mYCRo06MeSLT9rVjqFnB2AdnYS35AmC0Ce1QJkA9FedASu7B5dsdc0y26wIKhAxK
w9fmQQ7OrijZ4MzKC9saw6jvlXFCdeUXZODBzcYkt0V0Pgvt1EYoKCGmeT00ro/H
tr6xdFDHCacXYi5iJqcglo/WGchf+gjSzbHKAe8s5AZG6dfBATf1+7i6uSX4ePl1
cpJ2sQcJVbjYAxk0Vleamt0vRPoteZ0tAVJ48rmF9ftFivzcNxY8kLd7KMclEHOS
3w3w8AytzCvKJMclb8xNd1f+NLlbLevEkOiA4fRfYeX+aXWV9HDSQX+qLy5U/Ei3
wnaeSSrrSmopkKw1az0zGFrK3/0PukSEkInQhcRLDHzS2ox6cT6LGpjXcSoKj5nP
IzpJ7Bl04IIa/IDlOSqdqSRi5ME+DVVI2CppTz+auUTDpzFEZHDn1ad67I7fQ22A
lJ56iaqfkSjbKgAojhl0PAL5wauzbdbS0kxHDgTPuUZAZhN6MP4NzQXHHsLSwGyT
3NP11kQLzWreXV/VT6L2sXhfyqmGv1QKQ5w1bKFGWH4YeKQXFP/ufX1JsuaLOyYb
ZLs+3tDSXCU9TVi58303EiefZQVVse5ArknmcVOyludToM/M0mAg4EtL5qJlDR47
BhSHb2f+8gD8I9ZDWgN7nSDNMp1APgzo4Jmng279a/KlTBl4WgenEMrlBwX2X/vl
HxX0Qm+8vr9ua9xVVn2RqWMhcowM0OD9HRFqwuKKMddx4e+/GdBIy+VPARD8q9yP
+oy/nY0YFFYBx6tj689WwxX9jz3l38+efBSfR8JTi6SJEMMwGgNYf5qm8uqlwIw1
IJc/uz9AxNk2u4YDDGcjS2DscOBVQPiAZPdJjaECeKKO7bHaPS9ptTw/s7HrkEK4
RJdG6tOplrzNkMZJb6JUn8LA0DyLH+fUjfsbUq3XXAhrS4LU9djdOJR3gI68eHFF
IlsN79MvP0zg+JBx/+wVbVM1b04YUr+wQ3+bwkaIUcM8tnE08VUATsqgLEy8J+Wt
ic14DoUq78I/GUP6SqtpgO0IM3uozVpMdGyUW6CPOpNc73BnAXdGlt6Ujq8A0gX+
aqWhHqu9o7olYg4VDA5YmAc4qttpUczCA4MgtG2TfhIMbIbRIc3j4ucfAmU0Ofy2
mItPu2uAmCOP4ypYlP/UaMJX6PW3lr7GfxCRWXW9Pu+8oByiTTihoanIvMyGp0tN
8I9aJLyawGWfPPkJhaXkVt/GRjusjpa2ZfOvLpZkWQy2I5hZNK2RZ7NNkdeH56qh
EvawcLey0gtzQ6bhrLZDDd0U/MiT9ENYslzndaRBDkuxSNgMQfaDvMyw7hehybCV
s5LU9A4WSdjE2SoXUyJDnpYcbpVdSZaZ4O9AYMqAN75rMapGwYMNJMjz/P5XF3cl
0QTzWK/tAVg2mNR7DFdjiUkFj9+Mg47BGVLi9i2KTNvT9W8KIZhNXwMGiEm2qQ60
JF+ttrzDTOGWWPYcd6EEB8wtKZqIvjPerkYXHa9rlm3NzIywoUyfi9NfU/AJRxnR
ICXbCfUaX/38CtI1X8d9Pu1Gux2nD8Zs04qWczqb54dryqCYQnnFnc+d40YzTDwD
kIf22zSbxqTOzolOz81NQzNYRq+19wsIRN1He2h0o6BuaxVsYtkq8ua5phr1snJ6
h+62D1x87V+Vt9j05APxxqSc1EeOQfPtXuQTjz3doBE0LkGGOcXRwJH2jfS54htA
nCXmI0TnJUCxJNXeFU+czcCDaX3GKLX1MxWLyzFinXvJE9U2wS0C9d9HXcqBdJ5v
modfeRQWQBaJtG3sjYUoyKiiwpq4Qm2ZfZ1gh/ZI0t4gxX0+7mHN+MQQhEIT0lJc
ew9De74cIYrzc8odxvUUkbXMi6A/0ctSMMS3pJyqUxMmMzEYL6/NVIovIb+YmFYr
PFcqb+4/Yk1rkVjvdQKZwt7WJer3HAZiA+sj5JRqudCD/CyGR/KberIVccLudd/E
7xknPLZ7IQ847q7qQmhl5MDpDfLyjdIWMJrp8RkVbAtl/6jPLmyP6mr38ebrrs6W
Un/nifxx5pZYOxJMq2KVOmoELk2uLcLHbomH5ABnie9CrBlm0vtkI5DzQP9n+9O6
qUcDcm85eKzGGdf5NL2hu/jw4uM2/6QW87at00q9dSJ8mqpPWLKzdPTZ6zhz1Ux6
tS6/NXBCkf/gvCR3M+3c5hhKvjJvrllBS8L4IG25x6gNK9Ibhphye5gnB2957vnB
nWofLuJ2DG0Zzegnp9kNskwIqzMRjAhULkhBxzhehjG4D0ebc621aMgxzl8OHgRI
HjjVCfAkwAB9Yua9LnAow95zZd+06fVFg3BqCCQxEoKoRzjdXCEEDTDuWK4kPFTM
6SyeFptc5hZjF5XNSJDzJoAdKyHwpQsgi0AqiOfTf9iaf1daLv9MczoNdp82Oz3X
k2EXSyMvdtbVrp6sEZq7IrBKlI3tJ2BAtXjiN+53XzB8Dic+Khgs1ZRI6PSUfQit
8BzLjNdwXqd2l7R5DVMhyxZAWjCDUpmZ42V7MhCtXBPWx1wOSmtmKxHZYlSwkaF4
T4DaeMCA0et4buG5Y6xPChiw8zf1dwKpHZVs8AxNNMVu3hsG0RyUfv2o7pFSKbFF
YsPBcF2/ajVFHszTeXXCk0kAubwiCDf2hXFlF7qyfxg+urbrMBrmFl8EQ23mIpNi
ozbkRr8iJXj1ATU9++dV5KeGjRDnqnyRDhQkVmYCDuiqiv7cpd81gt91tBf/LJxg
lyw7F0wiJ3/hdcQ+DAE5mSxc5gQC9Y5JN9hlYg3SrJ3TxzuhQhiU1FcPxkPlqoPd
vYY148DWaIH1gYAQBnwqA3a9QHSYCJ+LNY7aQ8PgunppKNY0dKJ3Kuu8je1UjIqz
qZQjk/HNmN8MBp4Kc2zV/Bgl5BvDPAGMN2Ifn6Q9F+L7XKVWTUvlmc2Ssy2WpD/s
BmlSiemw9jrNfQCjElS+7mpRABckAclLD4dp9JvsMjow/eItUtG5pY12cbf3TxlX
85+Qh0a8SG9axIIIMWDxSG2Qz0KyY5gZMeO/lzI9To/LrdJobnCegtxKq3fu0UJ1
vOzuWqbsJylOeU8jGT1ouTPD3+3GoFePB0kx+GtbYI84mtyrVGMOfOBIPPYFK0If
DtKh5AX0HrhT/NCnLvoz1whSrSbVZXrbaQzJR4uamD01Spq3Wxkn9wvJpeZw+yfm
kjpDxSoHxW1NRTHzScs5bGv04H8xKIfOVGHkhDYAnsLLxO9WCwfY2/XaQAVzKMUX
DQHOMiFMWf9wROlz8ZqlV3atOub0CZlTkXIBI0zI9ZVH9tHdVIzoh+jbo6mkRHKb
6yq4BgI6cfEUk5mM4Wv5m9AcYdmOmPyLgFqPCbAmgs4qcpPRCiDqQiJ91yFfQqhp
Qe1EzXOrAj7fHDy0XIrwDmdEg6ZFS2eOMrdUYvV3Nxa2lMYOwA2fZ3xs1xOq9A2f
NRkrjYSLvHuKQwMUE7glUvKlYND3/yN4Yoc09KyOwtXQnhDf0yOhL6cwWZAcwVHe
M419INiIc3Rkqg+Afi+ya7J5z8vC4awsfh04sFXQYQGF3i5RVNSzRSDhkCwI17+/
i62XJ87+WjkinLcU1QlFNPpi2KA7Zm3N2iWl4mfDcnNlwek21xx/tlVHgv3dfNYU
RejYedijXAeA780DE8AfH+CeNXHwVOFLy9/2Nt4idTalPz1uy2Sq25byrY65Or0h
JJCrnKDy/hHtAEZ/yIvDYxKYhq6J8wHw0+dYPfyUSZeb58V3C2llWHtC/z+fvNC+
Gus6+tRjsyETzDWZ2tDp1JyN5A0Y/hiUK6vIErvjhM1oxwSzIaJggrd5QvUNre8Y
2i+qicA5Fa8p+4NRCnYmrMEwEl31lB/tlRnFuSfnmXTshdQAObuHBApVUIa1Mm+B
jxY6ipzv6L0m8fLEl7QL1aMo+3mdq68f0rnCE7sA8GB0Jjs7bc9iZfOeaU932Jos
4YcLq498tey9aJj6PSif8+konnjldbO230T8IduFiVbLGdkIxVC8Wp0mel/eZHXO
s+5WXyvHWTpyC372CAyT0DhETM5PnRfYaRqliKZoNOIyybUb/XnncNM5otB/gNkx
JPcprilzIH/pdl34VDDVmw71ks/ADC0+f1vz63oPhsZhz98FH8XmoBGe3BxDbXmb
CAEm/90I3d2nfogQLBunGSr5DgsM9N4ArSX96nYT+7rCQ2UseeZKWAW+1LHOqsOQ
3DeiSYfpc1jY8A/CqaIH4ZGuzKtUBakLMTektlTOUYoGY1Q3enc9MMgCThZkSqgC
Mf/g/uPsmmP9ucAvi2Xpf7BaC9RIlanrg0VXbW8Bwlh/TlUDUpDfOqkNo+yjbhuh
PWT9lqF+fRZUbk4iXgSAKFFxzrtp+FEbc9zz/3lzuq5VUYmEST6S9kTnWYHn+voF
0Suc8/dgyPpInSkfNluLm0IXClJu0iM/En2je9RguhHaiWnpq4LtW40j3mfeXg89
f275DuQO6JvfzuvkrSOswJ6A1o0zkKO/Wx7Oxrv/UAQu/HgYnbTKj/gU7C52BwH2
i5Ee7bh1B6W5kqnlb+EVo5BWdSg5wZQr2frCeXWAPxDNt5qz9HSWS/C8cMX/rwke
PBEux3q+dSwfVG/277xhQ8zk0PQxlT7sOZ2prsc7OnBLYqivwexvY3NXbUtdANUo
Mkioav1fGFXjXfQtXAC2+ZzapyC8viCLkXNW0hZdUwD7Ye7bYU1HPSeQMFfY6Fr7
c9RjbfBNzTl2ZOR34/vFE968XqDNqaMOQg9h2cOGz5owuElfdSXpH4mKyWrLjyAh
E48BdtsAqcf/2EmcCSpfGG0Zt7TAY9193G2K1xF+aITujIIb5xN3cbhAWFaB5PCa
Xzd2FG7CzVgujzxrh/GWEAYzeHcBbyUkbMAWIOCVM6wrMLmDqYZ//vT0ioFdB/yS
3ATgLUKY3cUoTpQfKekVjOsU0D/Tmc7alpPVrW+ZLHXpLARcFCT1A1iAd6UFYdzG
rv3Ku+0+KO8lcoIWgM6EPhGgqA7pkRQ6PPaJhfkM15woezcbjtPl4irM1Iy0T+F2
jA7qJw5eZM0qL+HpFZPJB5zr7fO4Y3LUxGMdNWlBy4PWubgxxArrmvUy+UEERQkh
UHrp42ehkPj9etMDtUMPxLrvjI4M12YZyKyKHzFf+Q2sXCPw4S06mGbmZPgxlfKc
tJeseVO2Sml7CvOPnSzIVDykg4SK46TzmKwD/10UVwa+laXvE1j7c3af/KEeavyD
fq27lBA9M5sashTaIP7Ucw6zlzyYTI19AJ06jveMF6yxM2C4r0CRWEEwznpwE4W5
BRTnvCUnW2ZD+KlXhZxPl0HqhDHp/1aONlO62dcKFuqFuVJhWXrs66xR7+t5JhZF
KLznldFFP9mJR3Nu2e8nKo9UD4ts7c76oFHO+U04CGyIloJymfA5o734cwHcNZoN
Q/JHIatSyxku9Zfolb28GK1XF78wA9iaN/thoMNaOOfWMp3JGdISTdvCmm3+g6MN
nHlmFp1PiZEOdbgq6t85fsw4TiSHHqShBDHUf838Zk0nMj7jnncLvm8hcap0qLqr
GaRrfxuGmaMwDBwI0a+2H6BQC9dW4knsEghAy9aWyjmDFG/TxXgGJjaW4Xo+sua2
jnS3Hlq3w2R3zFeykUM7/FdOpJF6KRt7Jdnre4mririZ+flwZwcu2mpzBVJfucy4
vPd23CRALPxyeMBZSO1C8N7fbQ79YPAAE94Kwav6QL6GeDGgjUx45fM9IOCw3omR
IgbTI7fEqlY9RgHG2kHeqjU8AI9Kjf5g3zTBwcIVJdAxLS7H1GqSAuxKC1UHJKrH
xBlHRV9dDGYhKVMR4yOM94gkLSYO0CnEpB81hn8GehO+abNMU31FQRggQEKV2C0E
zWuzmmGzsvpEV8nJUyrZBz7IVCM6ixlT8frin+7dLYsy8L4SRvgtcyAkovv5l8aW
IBby3tgsIq8fZBsSP7mXKcHn7BDmrykTSyhgo7ekFltNfGwbpWpby+b5mjTZwpC0
dmCQO2bXxnH86/Qz1jgAFEUGB1hJ02FmkXapOs6QQM65v7w6gE8L/lMNAwjtCIBw
O6jgzhRqsxp95EhChUy+5qGVUrJX5cuPXcU9hfaZx7bHqANhhUNW5xIblOFPx9l7
+1LuEPuvTeQRnI+r5ie8JezF/r9rqu9u1oup61YmCAk/aITG2f/IWaSjWNKsctsO
o1mdsPD9QnVqI4YIrQd63aiq9RCo+KCFzZJJ00cRO1ZMwciqLZkE7iHEq4ZQLH91
2wn32scS97Tlk4+L9mL9nWzwuNYHYQ5OZ+D15Kls97/hNJEetXLdNPIGrPzxoh6E
FVI8LYIOTBnKfiQYIFCIdN+335bV8R4TNSZXksJWWHEhDXRhT65SrF6X5srv2gQE
Di846QImmwIct2+cfsxNDkQ8qEo/YgQbt0On3om0Vws1Z4Xo22ud+8rVMIfKPBQU
UK92Nl4maQAxFARHLZlJqC4TcssJKYEi0ROllfRJEHfpsx6JGeaYM6qaLFmQGGYU
c0enqGycXmVGeRkWeQpNqsJbdkFvW2IxxkMMuanAV9da7eBbDw1Yxt0LAqryP6Fb
W/MAjuNLdIWMNVeo3CMp2bmSEW2tOGTQwNwAIiU9PLmxEQnls0zMpEBs6mIdIqtP
EJwjAlgsiN/r5GdnB7ooyBd5fkmBtCGPDAXePOWIu1FYoRQPjFvTTlhvp7XO+W7R
ZdGQpcJkl9QpguXFz6hUurK7ulRyjFikbCSz6Qn4F0aK5yt29/LK5XBCFp42B79z
FX0KE3rOMWQATBFcjl6pdlNiuSqkuwhibQGPFSj9DufrQEPL2Ee/AfcsI7txBJXr
SVVRL8iK7JjQ4ZwHQmqS3F6ynMZEQTAvBW8gLbXF1PH4vkSSeqgW0Mgp8w3AOMIy
Nhr0F33J0FQpHr/QXFQMs2pREaRzAU5NT1vpURHsSF4qmTEPjUOXeCTxhSihlcGR
CeuS/vvPztQMS+zbr6dYf1H27vKUxvVbqKWLnVgC0GSXAAflglL4Mm+b9t5wz04b
eSoNM6Ot/oJ8l1X/Cn/+c1yDCDUFQHG309QAlKxEwTJX3LvsnlIUkQND2HWEECzt
+oPFsiMObEx9/eDX37ERMKybyE1uxEWF/VEJgIypFLzCoWu6HEOJsW+ivQohJh7d
plf0UgWW4b9UTKfGcgA6uINs+W71T2zJ7CzNbWm0qMmpUf5MXKYOVJTUSzZX04Vp
DKkcjEhBUVgAlXtRQP7e8XeF4+pNtEHANPJ2ykl5f9rDp2V6j2BiLB/K6FZlwMNb
hPkwZX+yIRB+znmkmpWcqpUcmUm8Ffo+plRml4q8ENcFZahNh5LWcek/Tbrxye1X
62QBO7X8JY3inWAbfDE9vNKhDgZuUvwodhiTiDQ7KqX8Oa/ZZI142joe5cjrGbVM
okCm9RXnF7gUCw5SoRzdnqa1rR9OTtqniMUGqRmwvDItcLUFbTlCcPCK8bkZ5wEx
AMTfZXJ+ymzxmm6o/L8/w9TU+RTrZaEdZjyCbs1oElHugggRN594p9ygq1ZlxNIO
6wiiSSe1Wkw0bM7Bm+15V7S2kpo8ac6w8c/6yQqNh7GYx8kqHC9ZPRKRKZfjcuM0
nW8oqJad/nOE6G3EVDIHXyd5nHZLgxqYftMTEcTUTSwYFlf8rvBdzHB8ZeoxuNwv
/bW0e2ExWX9JFlvgxDyG1C7EtVO5DPxEmHjMFkeOZ+PvF/a12YgiSKtwbSEB3N8D
lHKfcvIj0x3mG0b+w3zmx0FBpVMVs2wVZakaJuDjRlVM8uZIk+D1p9Iox+FkB+m9
OnNWjeSdDCIOx6B5oSc8bgs1O15EJ0GYf+MlWOyY2jdw5XbtnyXQEsVE/AXvevOo
h2gj5tgqt3gh1x/OTma8wdznuHJhI0/D8/ykUmiW7aoyBuQhW6udBQpbXFAXWzTZ
a0QHFP7TUQ2zBsdFrx30cWmJXNUD8RRKLMiNFX256c2tL0GF4hlOaxvWIM27tGbt
18nNrcE0vWTYXjze/Dzlwwk6en4tK8oS6EolKqghfm0xCNa/7Nv3cwosuVZGPG8d
bpeRRpeMtiI7hcNFzZcuB545tMpph6Ak1RMOcV1AgwuD56SGHcpvV7x80yJJ4jzw
H9KAIkH+mYA+3iVvUlAZpoovdq6fJEjv5QiVujtAAFh4Uv19iSVbfcAyDxabhZ3Y
zJm1jvHR212OqfxLOnFcPdKljTe3OdadbxXjjkfstZui5cKHUuq+Hu9TgrGMnZj9
4K8iLs5kScnn4BKrrXSRGE3lP9r/J5cPsJX6z6gxmmPXJxQLNSm+afL3X/19wAOV
VgwxZKXpZXoHOfCCpcOrnxA0pBJA5/3zChU+/MgT5Lt4579IdwQUY+4/rPtHaoAs
xHluGvAqOJqyydTaIWFeuxwVSDlJby+WAVESauvvh/+YssYUOaFF/n77fMem8NhD
G9/ZLPiytQ0F2sqGaFP108CS93JNvjCl3QZm6TRylujrHqM4MppOpM3evZ4cSnGu
1NJtQcgw1C0F3cRm3wxLxZFfwQIw7rL7MgjMrOZ8S3cZHImd6Qqmh6fE3wCpnieu
uJkbU/ZkOUvHWoT3iP6g59+brZFcOImJHT46kEMeJegVFH4xWoHEZqeBgC/xK7w2
Ju8OREd/Zxmp6mCnX2zxT6mgjXrFJSuwkMpYp5IOMusApTYuw10pE1LMNJfyoKTj
CkQ87b1QjmQoMLUHjhtzfDEGiuMgqLJdmF1zr5iY07oeL9JoXGsehJOZESQjqBng
bkScP4RgT/CE+ON6xUaKZf6D3Qqt6JrqomgKAwfZFu1mF+6qjEShGz32FvsoibTf
ZDAo6BP7dvX83ah2qOssoI2G+eioDTIkVhKXbFmYt6tuDFqZzMjmN0C7xbwaz77b
ZQDitFQfBkHMz/6ptiYACEv9dqnclpzRvqsvQrtyv4FlkP0KFSmMLQ5XIvfMVXg5
q7DYUm6leHCxhGvMFYQVTXLDZWdQefDa5MFnwj5Qh2v8jEABwFAfAoPukvhjCj3R
RIUXipA2B8hzFOx3IV7oJqfO8BUbt/juWCgb8hIWWPcDGBQVpgZWsG37m7sx1UGx
8CYFzJCE2mM4IIOE1RkVAftz7csUVnXhzCD8UwrhA2EdTnB0NmNjIvnNcAP2J9fM
JNiIS6/LXrRIl3vTgFuhE54P3DbXQiWXQy5oGYxCremSZ3JBsgGthXeit+64X8eM
LwN5zgL0P2TqFnFxKrjYtXwxVEYo5qEJXahILGkiMjO4pqMA+X+96CQ3b3iTo9Bv
GeFvNEckP6CpSFzVm/t7pxIKOOu8GHOtkY2Rg+k6GkxPR7s3sbm/tenk60uqSG+a
TwHjfxA9eFieAhoIHEEwMvXU7z9+R0NRQjw6vopIIy5OGa64Vm4xfAlILVB25U/l
EQxhbyVZGKfXvkgqO65lO/AIAv1KIRS1bVtl5k8fep7IJlmHhcqYSjLC+1HPUkbx
pXubW9zTBDRUuILGK0/9kskmwIQPoJvg3u4iAIyK9Vvl0jHrTO6j6qXnxXq5thGg
elnNAmjeWfOKHsudpLoViG2Ob4rk8QtfHh/a8GsaI6dmvU53RZpv+YA79ySU2AUd
Uoz3wu5dta9Q+FHXCwScHAGcbM2RkaxE90OkQUhBkFSUcEAMPOPAUZlryM94okSK
J4wcAFAe8RSf0qPLYIwDyZX82n9wxh/9TOMAYGADIEMKdBEV+6/2rFGAFYC7o41R
WAmVHmnLBSCwQDc84y4q7SbAgCYqrHo0SLoPBZFEgEAqtq4fdOJ6P33u6o2sY31b
BRrJePYFy1kBnkCsEMfcLWql/thZlFYZbM6AZ6ytC0RXmVLLNSEkU0T9z9jM2jnF
zdHRTZ6unWvGxPZmvnwMoMtTIKHYzFujPi1bEZ5g2ZFTD675Ob0J6yO0/74Vcuuh
edXBAr+7SyxgJG6VKSvwjKhc1nNrCZIBuNI2CwdP0+6cnywD1b6TpyldEMGWUY3U
c0OGAGz0Bu8ZcklSntrD1CEw2wIUGnr46CoUnZTbLszmcYiO7E1Ok32KcNXwxEAd
u379Cw0O6XtIYv5sFUPnlnetMSCLU1o4yPCxpMqPcoMNa9RgqwIEguKjP3wg51/v
8l5+IT4U73F7+RVyLzhCjZdBaft/Sx6WBODbALYv/UkR4yz+6jx7xAXrMXeh7x5X
iZbnWWAzSsBPGqfXVfds7rnVBlSWt66S2Jy8TEc/RsAZiAoFcB6pBmL7tP1Mn7Pf
kPHOJCSJCcehJrl4Ccs/M+BFk53ejK+zRo91tiRqorWw3wwKepAuTkIzWA94jzqm
hI56qEIU7fXkkhCIIwPYmNvee0hFY3hmxk5LGcr579ZyHWoIeRDf+GfL6P2j4apM
akpnCQpQ/EZ5Kn15/l7S2Si5FqupGra8XT53y1wPO8YzdVuK7Kl+XxK1ya3MPL2k
ag+OTkt7mfBOJSLGKp2EYopQFL9pdV1VBMyFTkFjnd1zm77iC/m/x03BdeeSsO6s
i4+pSiHesjwS78br3L1Zpwc9sCJAX1ydhiqs7c+oDMj5cnfd5/6aUUoMEZ8xtqE5
K0FzH43uu3vRVYhNAVA3egTEHQ8I0mYuTgpayNQbNWTZ1N3CtdRT0RbSnev9+7tq
gv8LdJVWYmalW9gMfp7hu8/+YWjevCFQGbpXYTv2F2UvQfnEEYaQNadOmgG3SXTC
Sb3t1EF1JEkWPeq3p93wKGncTqEaDwBPyyErkwUDxX2CnXyjT6C3rV0fCawUJ+vb
bKijRTz9TGYfH81Gl5zzokHy6Tj7PStS9omP45wZ/iu86t2BGwl4gK6iynni7cJL
dl7slCpYXJAJBbKX3ccYF+8QucmqR6mlUKdemfaExdVwnqnqRA24wCb+n9SVzEc1
54mm4xR42KyHmcPhApcNecHV2bviSg7g40tOAww3VZJS1W8zDoRggplMnQ8WLHVK
rBp1Y7fOd/hdYf1ke2eE5N57w0TKIlkYBUpEA/GBvUdM1SOb6NxJNeX00dlXdJbu
T+T4TaizpCsIYzP4agRCaNhg6NbIJtbcKy8q4Xy4HwNI7Z7fEwKF4LH4NXxN4EnR
TWgYbItzj/hVLsioKZ7AzJ1d5nCgPyENkp4MbWJpQJx1hxpV9uv6tXrFDHPqTQWK
isppdArWh8HtAWVf48dFS9p/mo56rCQvvqImRrMDjKFhgvtT32Bp0V6RxBvFlxEy
oOd2B1bgdVGNx4pXQs/nauCAIYWHA0vgobf5x7bF6c6q/VHsDOhGdMY15XDYxkSz
NZFPlkNT3MDUMv4GKZ5dM0zVtgZ9MXSx6ZJOxqqGxi6jjX0SBtZ1v4bEtKjXs5Lo
cnMs9jdSQS70j9I8818sNKg/pO9eSS91XZBAJHoJ2ScD+aLe0DMPvWnMxBhu+RgZ
9wd5J7os48PzwkNrTUi02vELEtmRQr4bJooGAAQZhsA9i9VdBBza0uchSJmuCFTt
dVdS0bbtpBectxEjOD7iDnBVF+vkquyHSzxsmJfRLY2I9WZwWBGK9sC0htlKAWVw
8J3EHiqpfRbe29uQgQe3eN0++CODZkP9QjxKi4Jce9cNW4gJZev1H5gLe/fxzeJG
d0dzt+ggfHBT7iUZiU79G3QyqksEnJPXHH6vOQC7qlXzTruAeGGevtjNNq/TA6l5
59+9KZsJxOcXRtWc8UAOgKTj3dS2mtcPr9BItokK33wTVdVo/18uFcicY/x6HjMm
UbeS64HoId1CfRAQz7htXobfpFG+g2mpevsNaU9HpHV4lCRuVH/I80HkilbOEfXG
COuwCOwAlVYabjCZuwjYcZIOfI8XAJ4H3S1h+S8z54/uEBRJM7fggy9jtzW+y/MB
IQjWt00RWaw4cT6e6ZLuzuTiEUuypnCsmGpA8nDHc4MjI0ECdUtn6gDszYLYgaFa
5Fo0T3D/d6L57H9zX38O41VoBsi3jpZoIHzU5+Z1mJRRa5w9UlMXSG3pUU1enARE
0jpp2VulfW0BE3z0YIjtKIgFvGQZi8Lc3tq4TAi6fk1dFpLPzCMAbWnUUfTg9UQY
ZwA37m2idYfdeef/pcgRaGhc7GrwQlMX5ah8dnBHz+1Lw2On0fL9twTMfxp+jKnQ
/GDn8epU7s5W7lc0PcNgbjDBpNpG/rxrgvv/3IninqNwG4cA4QqdgQsPiTpFRhgH
j5bJAgl+45D0l+KSkmfL3hf27r1RJnW9qs+C/i2wcvZ7B3IZ9LhBIcDg5jVYnlGg
gqQiM57jlWK9xP4lJ7c4C0HXaE8G5HPeUAPAubOCOMQC2Yk06Hr4vH8tW31+rVvT
9mqxk4zflmkaAGERmeVMDhvklppBwIJVKjCeSe7qeufhuUUr+vpLU8Z9Iq45QcXA
Y7d018rSuiyXD6CAL4lzMdaxlgORyNEXyr8FnB8F259T/riCf5C2sO1/BFB6aj/4
ObG3/23M+/Zo56HqTYVVpw7WojsfX1fkyAEDCTREAis7rPSTar+q8KaArFu3GLwx
/2uyok1PwiOzGh4WOD3tAeGdLeMCZKV49zAQv1eCgCEygTsil0TufcFoWJ4/J9Ak
A7prStsDK44I2RM8cl2TaeU4U5yW6NyilgcHa0SwmUhTTQyxEJwUxUdNn5Jen/B0
bTl57R1jxVqUfrOPFMIOm1DvGMS9ucFxGKRhYPTfOYizaNgD73X7xGZeLAekS7i1
KSsyarjufxC+ocXAacZJgy6Ar7Ev3SJ/BOVsNzdNXvBxcGNmM9qhoiZTXGogUPHt
i3n8Q0KVaJ255KOx7qyj/NpcRRHESN81GpSIB+DRiqs3sH7cAJHDJKJPhWryE/mP
docgEjUDfkMMJDgI7fsHTj/vVYg/+eDJiy5APg0QuqFi4jsObyl/L9D6Gsd7itVO
FJHxI/MnPR2wJAG4XcvoXUtIU2nHK7lE116bb6v2KfXVScNEY7cPaS6KHRna2JiX
8fuulOgV7fHJlTJgmU70BU5fVNwirFX7f6efW2rdvIOfskjGvz2Oih45mlbFBTUz
a/pYdQsgEuTNnVH5ltXNpFxWy/tdhH8D0t8+lLrHp/rf4dMfAXO9fQDy9BYWI/OD
UbVv2AlFlqJcUxR3ibhhAWFTykrLkAKKZTrBY97E8Sm2LYISWuD9kURHwHsAb4Tv
RMmxYAbIR8Kec0qRatzlLrTwqb4YSCZZ0NwQrm9ugxg+S6tTbpQZPVjkszUlSe+i
HpLlZ2EQlXmEf2Ro/29UmUITrrKwEo+SzsAsTCrpiy0g/ynzSsnbkBup0h6RnbMP
NYyrqFrgYHoqShOXLnYGPlbzNxmeaZvFjohtmNm0oP7VAPB7gjZY0CSB1kx2w8OL
aHbA86BDXjL/k0Apir4+sSF2flOpOeacYiulae6ZgY+nLavuNEQ6/RvetKizqSeq
oylD/3aASRwyboJkJUxomJVWdZJvbrWrZtapayMyELR7hHf6aAakh2r3hPsQjRTo
cexN2HyfXeHLVmOLT6Jo+VrGAiZOtsoHFZ0XgGZcjjM9eurov8GHKUrfNvadyuTz
jMZ1VsXecyDCs4A4S6xHXQmvxAciAWl4M9lS3krXdHYlpWqE8msfWbJtXMwp3liM
gOWGAEMre1LHZ27X2rAoaN4A5TyGLJ2cFLLGh9tsXCHMbRsSw2MND4wnBM2vQ4OA
MW6vbSsVbzfKxfCvSe2yi2/jFgomHk1bBInxoNAJW/2slpRkij48Qy5yiFnsAOiu
d5wu8jVNTL3QmdNpd660BFlaUyKLxB7Gem4ocFiK4UUtemF870mh5CTsq5w4Vwln
7KymczY9ayAqr2zCvrya2h/eclpnk8732J5L1Rt78kri4HJlkvSH/czJg5csSGYU
1iobINXMSLp14CpiiKuO4pf+MyzzXjzGzDqTpmUqqpyYMQaZz4VGqMEOMir6vi/Y
3TlLKVBdx8kqDOmeagOyeakwf4l0yTB5wvKve3dCm2cfdkTF5TPpxsajDCAywx1a
R2yCdBdQZYEuxusfW0W435rBwzyQK1dUGwP8RYBvjevJZFXhhnkkRv/9Sr4nldFR
Icxo087hVybH5qBzkXx5RnS9Y9XQVLClpIlwyxlK+dSyzKrIC6xo2gATrKbL/HO7
/rBi0YxdSyn88iBDYo4K8B6GCl7xwe6MCn5xi4kjuJJA30onbPi9w/zrJbbfh0OO
MzBnCc4V2IGR5deYasqihymLYFNSIQQVgKoaKbtuDyLjm9zW7aJMwl0ZE2PFwbP7
l37u2KaqiuDr3JZIbIvwoqHLY832Taj+E+wJTIRKe04L5sK3Dt4jhT5SbhZ9pKIb
0dIIbNgm8V/pqQogGRG0bfNpTXeGD94pd9LZv89FBgyOzHYFmGsmxYigJFJ1dIvZ
pL4kPJNd/3NbMMc4mK53IkAENkUyC4p1GB3XryGlvRsBeeAabmrAU0XPZB53++XL
FoqukGgglOHsAHe1CEpY9Kc7zDg22Ivrr+UvuqwNRMPYLxmNKtM1reWquCOzMUFX
7ZP2PhbI6AFtRcWmYzEJkwBdQTCs8FvfLjb7kDSM++/470SLz+WnvGc0qIV3EBhg
T5HFbhfB8wWXXdcwdCePyE6/7Q/P1QBAv2k8odm09hbD8TyEBL5EJ4ZRRRIQHdao
p6zW2Atw3nO/uB6M1EBUw+gLQtcT2bbbQRWp9X8SndN9SXRL4Jm1t/dRKj0rsCPU
zjnWGfSN5F75M4u6fmxvnWfCSB1KIj3lGN8DX0oR/m3OeMyVYQDU/GglTPIm9DKL
Py45i70Ez4nWXJgtz/bfvnvghrR9Xm7YNwH+pZk+SddB86yrBkcl+7UYyYTNTmG8
0NdbNu/LfRIu9WmapQF6/zAAyH7Ao0AO8vDuzz39dYtThKFgwQcPqZkl2oaAaHsm
I4cApKiZOBwq99WSIasrd68RAVQNSOeUkmD4ObcslaqOl1wW4PTkbRkydB0FZvqE
frHDZJPrKZ97xnqiHv3FclW8dVxfI1ttVjNfvy0vFJEo5trGGmcxM86QjwW49kdW
cXSdJMxcyPPDjOOYLoRG7B/oK/dVIk3WatRdbY3C29GDpvCo/ZFuiuSHjrh9jnyS
smg7AkG9P0fXSTgIag488JEo+H1WVjhEpK85GGp+uzgkpVniycBvN8raibh1hath
82fXMMkpjfVg8NYgf+DnJw3wIcHtiwt/jPnFMSuog5Xo3o+hJgO3yrMARt1MCMMG
5evNsiXaiNoK3g7dXFL8OzKD5IrFQ8+/hS6IaZEDcos5cmZDYg+GW6P3OcnJi3Ai
dfxwRnS+dqgYno/4rc5fbsN0N7/Lw/i0qBriryMbAaLTXYmnkjyL7Rdnwbg6IHFD
jpsuHT+hXowTh7DIAayqXkul5hxz23jjyknBoWR60yRpX7mRhqWrD43H5A9d8OYC
sgSblWahEoMaZJvlZllmsaCCFA9WewHmtnVXCXHGgsCBx8EwcAAMFEIFn7Fc8d1Z
bgVg8zVEQDDbzCYBsukSpmaqQBHJfQF+syPkuTneyXyq6JEJime1tA8yU8G1OXjw
KY6Lsr0nHe8rssqNcsurhpdKIqLEW7aARhn5QHT6AnDeBwSPw3qbOMF0HkpagEo4
CAXC0pmjphc4pMUo4S3SawdMRw6551hI74Q+yx9b+RYyhiV3nd4AsaIOQjo5HIeW
2njrud2e1XdaKQJBKroEA+gtjqNto3xDxr0OlP6NdmecXBr8vIht98CNC2FKZcvt
TaaASxR8ofTZ5Q29lr1KFmodFqD86GhNsx7CMPoYxRC2hfmQdfypCbvDiC2rRNy0
t1DrYLA8VvRF4mClXz0IdLfh+bb7N2tybyT7DGT7oSdEUuDooBTaqryc/++RIpB8
uadfk3tig6tvo47k2CjTPiGbXw3LxEhC5qFsQmxzBGAYwr0Ida7FWR6znEfHmDYb
I4kP63CfnBXz8uAvJsa/sGsUkJXWizK/B9uFKm2YT6trcYYmr0cDU/HB70+cdOGM
Jhr9k8Yc/CAyFzpKHHpEja9zIwrKP5fyKdNQ4/O2Q3ZrOB6jccUSSTjQ7wHHRjvr
wwsuFA6XYuouSrwJKOZp+G59Jps5TBpoIfH8gsPuxVrAybdu2BSGPMhgkosHtQfZ
Bcn91hBOptHxaABiOWJasjLYJfJUDu+ozOPW8eqDsSJgW10hsarBy31Zk9MpnKB/
dKJ+jj9CGOMGUpMeBNdCONhaf70xrQ4YIBgsq4UUGp4gkrHzOSmFgwxoH/UjdPCM
m6qWsm2Oll5fHjFeOh74Yp+WSOytvF8AI4/mtISiOas0fRe2YUFysh6xFWBOwF1G
IXKktwUkuaQESPZVAFXFm8MqcwIIaK8ZveEtiA5+bBXRcJko2wX4aW26+ivOPDWr
TuXVi0x5orVyTFT5mmsJJpYdAaQJMo4yMXxQqsjUf/XSjnJX3wW0QskP3xGX2c8G
lNa/zCn2gTazErzu/IKPg9+0JKiA/KsLPoZLhVguXXjoRRlpWnZTSXsVpu8GfGnH
l1Z9DQ3mcVimvK4RaD8Lxi3Nfe+huwXfSB+xAsEJ+Ve1dEjarIvt4earMqpRHllq
pwYrKpjs69kFVmf+tmGcWTbRSMu336/n1Vjx1mCLeOE/bDW2n4zCH1i7dXWqkH3O
pl/ms6PzdUpjmBNRPD4AX/PhNCk93Ql7P3oYQAaNhRTLCnEwqLLOQxoWJg2XssRh
tgaqmUIgTzcsY/VTcIXfF8ylXQ/ieQAoxyGRkQTVvOqGUVronaBmEy1NIVstenZx
HyTiiZkMfTZ3NbU9qKN1SRRSi3ybukEKnnIEBAmBymLl/AGfvLkeYy3LIxtrzONA
GEnQPhkcAEUNCXq5GZ6/SGQA9+Jobp+MihHWcYIL0fJ1GDptvvbfJ4urQ8zRmkjR
/p+l1nZ/akyqCKuVoCeP52VowxlWhBSKjNjJLFfvwA2zMXaFZVae/WgsFSDnt1KT
/MCzLfJtSo6Cbs12f+7cSGRYNDHd7kOXwMnYLhUnjKb3BQQ6TIsODPgHFPYaLmib
6KUuslb8rV0Hc5vqF4EzLrQDhTPhE39klt3eWHDUVfWYhUPaXLbi380AMRGaNSgY
eYtbfkPf3knn6rTmeRz6VnjTeZeLWnQZpk8IZHBP0FnpuV7sDJyXl7AxYKAZPOau
Uox5zZp9DOh76+L5KpknlxZoKY/eiSwud7adUPFYDu+fiYoXVYi4Zqo2JKpUZ/bZ
peSiSZ4iJLw+Xgpwv+xzkqpe+5SJDBZx73JSOKE0RnEadIsO00nTG4s0yoa7Cpgs
WiefNwF4UPY3DGjh1PWiXQdl+IZN1J6roByc+ABbmWtdmJGob6SwAQLtbIb9XE4F
lrUQwdcXVAMMV4xz5Cm8dUzW0Y/YMbiiXCpD4meCdMFKa5a/geLve+FU5aBsTau8
4V+0kaklptr/LiVo9n0vZ9UCVWN4ZzOaTuRRxWsSYRwwYVupJr18qDpAXovwFdUe
FY+DbTfqtMRv5VTpLhRMtBmBHPy9TSiIpI/d8knQYg/DyI65mDYnnBHalZv9yu2K
PwwL7KnCWRCMqDBMHiaDnNHBLGS7ewOxwK+ynkWWcwQad7XOxdoV9M0CtxHA4uFo
fnRovuv32IlSfvg6OAMibm3ATllE0t+zl2URworFKa6DGbxTc3rl9gYqh60cooZN
Q1A8mdlwTGS0OZN/djdlcm1fbjqo+IGi+8TOsVUDAXhxK+GTmnHisQi01GmVgBZZ
plWFZUhRcoGV5txg29yT8L6wdbrrL/sv1PLGUrGyyf534bPGHyPhGG59pnB+eZI+
SyRMGDCYbFs5oJvnIg/9ipiIC1W+sQOsdDyRRgEM3QuOQD5Qy1S5I14bOC1H1rwn
+X8aVUoPwbYhxJEJe4YxT3eQ/qOMxL3OiqQtMlWx+UQl6Vp0I8aUBIj/yfbfDqbs
IRS9V//fGl/EOJelhgTBSbzY9lkIQNxoR10pnbmu8Z2rbeuKiy2J5zcHPHxCxga0
rvOAfO50LzmoqlkbejyLbsfF9gqCS2hjVdvAAngTqgJHrxDP+nCiHpU0dUMekqJ9
yQA4g3Uaxw+YlQt2Xs7rc6MPQReEFQ5mm+CTLBd44qBDcHiX47g/kYtqK7WDuLRy
afxzYWRAEVNIRrkY9uO+pvr5u24ExvGHc9emEL/HBu40RQGXgiJJgeugSgkk7ivC
TYbTmuINVgcGZuXMdrHqJnZBvPUCiZV58sk2/G5dYp6Byz0mGwdzvK7Mpj01hCIG
VivX/HEtRAoAyAFP5rpq5V8NyKY1PkdJACV2/gUaxt1lJ73UvXvv7gRw+Bo1oQl8
jv4uy+NAP7BDJx8MPUFKyvN7gcgtvfSpikj5iR5rkd/i9GBaRvFejnukEafj0zXf
EAixLSMPFpy98ECQAAWLghAULESdwOXRnQor/cZdY0ALt0sGeQYwAB6cUj6bQ+Wp
dBH8cBI8hxHJF9AQ0vXZc0kWhxp6bAiZ75MsB1UeojoT5JIOMbYeU8gltVvKtPy/
82gkS+76RxlQfHEgz0AS1qhmkGNfF0LOQTjDV42Qe+PH0IALKTKYrIai9Pox1mQj
GG9QQx8POwoxf1h5LmGFO82gdkXFxltnHwAQTkRR0z3/2M+xARQTi5PR5jkKhlYX
Tce05V23LnsD3OjP3mXIBSUkhfCobFr2le1s3XQb7SxYWXzksbmkz1bPthfgiysd
rvJgDFodOumGwwYRBMCX+noe8k/ndTAVC2LJxZCV+umLb/Bt7nrd1yRLX+R1GUlj
LWnmQcLuGBDpNtXtwBfhKZGQuf9raFEuOuewIrJqOXQH9Tr0jcYYTCKDwU1w2GFv
qle2kOW2p5Bthu1pz1xTrHzadCc41zpbKrYy8fn2WiNJEWurKvbix1olKSz/llST
pvnsplsgWRVTeFZBskHXB6fBZ+oFLNNOlAWf3MI/OiRbm0sNFOi0v/b+Qmewz5P1
z4+wg2LSuTI7QoYQN4ZIDAvVD0zqV2SOkUrRsI1N2OnzawbZeJb8oakew+dQP3tC
fBdzGZOkAa06mQaX+brirSxC6Jugls2pcdgd9WZ8KBZ6GdCiMa3PxdXhg4XXwkqg
pB8ikbSvpw7qUvvq8+UxtnpFDU8/qW+xk3/1V/0KFgP4YXJd7HwNvm9J2qQG+3+t
9wodU2qyj6c5Zt3R4tHVQSGI2C9pc9Fgwhu6fhQIdaGaYloovvNn0Bc6MBZFi1Qa
dxxDQNga4WIj3zBky0qxMZDhvI7TTWIY2F+Fr0iy3UzPIL75Zb7hcC+ppfNkEkfO
WKsI/wNx+IiDjrFvmNCOhHC/dbAMDbu3+ZUFmV4B7K4ugWTUmQGzYnWORbAfx0L6
mi41I4ZPYgJBWvujF4U2HhqIoS9ET70xdy3s5er3RpTZ+JAT9iBTY4X2s3HTVulf
5pArYMyKHVfWjz/1Kh20taFGglvn47SUPcFEHnM725NvGrf54FiuxxdobPS9c+nF
uorcEHXwM+vmdpXY2t8l/tfqL+fa4vedpWd4wVz/LE4ArhSf9Aed9KVZqfquX4FX
7kYgOh4+nmu3JBhpamEi22fQMwMWYkbz5Sdg5uCSpTTSomy/AEIMuoSwvLXd2SNP
+5vil1OPQjc/cKVaGu6kSSsTbHdsue5ppRBZL3yXEYu1cy1iKTzfaGJymkrLQrX0
Zyt7rLSFK32kuhYPeAqAx17ZZ2ffT/7a8tdW5kK1ls5nCNq/1z6ddymomqRspI9s
liMiw9dEB75d+PTUicfpVKRbAs+mAKJaZmDjH+fy8AEhjPYhsiQvu83bFBxNVqbz
vxCPwm3hSpDs74J8C6CAZFJ/Udsa8xUs7TpDooMWGPSl9aq2xBYXadposi9rAH4M
iNomporylnAZbi1Yoh0WZ296XsMQFJSMxtVfp3hkGD/nPcqPPjvOdG99UAYN2WcH
IXb5zYOtsdqo0paAXUcE7IUOBFUzHZyqSAV7TxQuMAi2tduruIhEu+LmiN1cVcwM
a2rLNm6FTSkXML/nqa2Tgx+wnOItyhN73luup6hCVNsRMZe4ZzOqQp3lgThLBAxQ
Awd3+5bxjYuloyhOY6VeINkCvqjPwSnYq7rdAFbLzgCto9izHTACntpGqqFUe3O0
E7a6Ol1pHXdCkdGftDcmCwuPuT5MximUOupZtA6n+twFJfZBmXx57VGv3iwW8Hv8
Xh2qTUjWpgvPmKAUrugo+bZ4vtQaX+R2QCaQDMhgB+FQpxicLNCLbA98kSuVCyG+
+OGBESPUjgfVzgfdnhew0Po5qK8sMx46kHTB0IYzn1V2EztiWVTWfdOycyGl8Zhl
9Jws4p+u2cKeGxcVQ6zKLDh2txIja2BTRebLFVWBo9/KAor7imxJp7kOo5J+UT9j
DSgtGoO/UKscHec1BrN4pwvhSYa0PVK/8yxxpVJnppm87L7DeWYMQpJIP2WvMH++
+6HliPXEe8GOu2p4DQwvhPxkRSng849zbsfyMJlAG5bqfdXeCiUg6mx7hXskRK+w
uY/IeC08GM5frrehaKr/VCwyfHFemoTiUGPwJSq4PgJ5ZUGNXILE3JdGRjmv2rp+
+FENcMaACRJlWUFBqeU6IClD54a6SYIdR6bI8DJQItCUz9r6JBwH0pGcL5nHYJ7Y
JZPC6ajEZf0AZaLgq/7j80Akc+FfDQsE3icu0u4DQiLhvQ35t8JZFGWXLV/lEC4t
9btEvSOsXj44sqr+6wFkoPGAYsJauxiLWHd9IFaOPtUFJDAkhFHDC9EgmdQ1cmAp
9Ogo5/Zdl1/srfZ4HihIuvMxYjr5RZIVp5/kDlYrGup9EFOmUkdd97TBks2dgl75
WpZyiGV3k8veTlRLE9XeTuCLAz7U1sghSDN31vuqPM3rk28wAo0X4tTxdAovNEBq
j62MFzcILcRxUe2VehLwyegGBsCSmZAcDIqqHUjLYEBMc/TqqJ4s1My2WIdh4Ysa
OMqHCoRWosS5CV6FGWPfL7dOfbB2t7o3reS10BMAyLJiVsFqBEuy9GRUkJI0Zv6K
fuTf22Z8XAF2Lo6kDSsW7Go/R1jzY5r/NeLZyIsdoe7uc6bnXTyLSgpPg7ciGC9K
0HTYruRCIhGWTBWpGGlg5j6b+q3mo5cWRrNmKIgQrtUaD+eRilvF5ru+FAYYJgKn
UOchu5XOgxTZL/84qwiPLScft7pvsml3wS5y7+m8Vu0nK8995bXRYDSBQ5SMDQTR
brhOpwRzdkq+FkLFTo+L4DS80eU76uE3jNehu40v4raHuSdqa8YQ/bMJOCsGE3gU
tr8OCoHnd6MT8DBWi8kHuqj6TrDF5+dGjsaSlJDzAtnb7fLx/6GMirEClLHB1ko7
E6lbu+u9edpixrPVvs6r1GxYpmRsuGf47QntAzJFLp/OUF0iO0v5DpfkzQoiydOR
k2G0cYykFoC2fMZmPi38d6CYNFVFXHhO8YHJWEr2TFkzYko4xlgUh0NvzZfEKuLM
IsoHdYRT6dNJ6aaaZjzFULqsfN/TdJigotWc+04fjveTxwlP86aA6w6sibMzS/SH
JL+e2lrdb5kE3AEfaBdlu7rUvyVSXZt8Qbw7LDiBFOITmeNCuvi12vMPx1iEDQvl
kUqy8n2SEozEYmZp8BHw1AAaJ7ULVNEfkLw33LiEUUCDS4z/TZ4xCN4lXkPigmyS
3UfLr5cxChLpe4fs5fDTHI5Tr38yyXXwSWjObf/Bf0gmMq9MmviebSM3Q3UveEy4
Fksr0rGsPVtfMF/GaAVSIVr8Yc6dZzh0Nti8uO6/UgxNn/Hngfuy+ZDqZVFoUC/W
VTHuEYg/gJAxryiabpIAf4gfGHvKpY7/MH5rXTOUZaF+F1KP4KzsxtUm5cxeERSU
wgFv/nva4E3lVShh1Mm8CMazdjXGwP/sR7MBM4PcyjExHftZ917OvE3DmN6oNLTy
W8ROK6MLxxEhh0CPAzm2sMcaBt/vmFBmaSeCWmY5e5Qc2IZq8BGp1k5FEz6NDQTq
pQHDG/b0eMC0XHuOQeSWermvQaJhCOamnMXxAvi7sBPlvRBZJr6mW6xcb2eR7umq
5ZB8GSLxJ+7xnwNoPOrIPnsiMeIU5wOPBwyRKZNtIxPYcHMCFhlNOLoy7a1Rgeu7
Z014h/k81wKivv4j8pCrcpMg+nVMEK7yexIJpASQ4Sd11eZdX63IPfl1mCYwbID5
6qzGVj5MHCtVTUm7I0tPf9+fsTViCaijJrsVAvzC33Sx9gau7OF0YbP2BTA6Xpi+
jfiikSYpRJEgBp8mbFK9Vk1speFANVzhoEYsQcYnAdkzWdXrepn/Lz0Fd7x8PakY
9OQ1NKHEUV+TCR58ELjUSRbMSXgJg8w+yvLovgkEFcvZPA+dg8xEXuxGWZ07k/HE
oRZe5jic0i28BkIxUv/787g/68ivu0jy0m0KEpLHItoWvZBfTZkbfWHWGaFaO5mW
fAKWo039CXw8jKqidLNGkXl5Pz4KsY9HS/kx50Tut58UwePzSdSnoyjskXl3shn0
U5Bw1027QLAW+mL2klfbLR5HrdotmKimP+zu2PkADZwbnUM48FGDvn2OoTuEA5WR
RN+EbKL2nwsMvCKRZIsudPRDetVxkHxsHEqMdytoMaEhgbiUtt+lVSQ3mwT6fcWY
7q+kdzSipvO4jBluJLiC8EigF70j1zmGvtlD0p+akMi3IChSguN8XRrb7YDUFUUp
ELMsusdC94aQ+6aG9nRsuLDBkQgAagkWAF94K0DVScFlVto2w+rFTV9L//p8119H
VJR/XTg2SMxHiYS6pn1cXqNP95MJT7hHgajMY39TYG07t40OrZXxolQPjtYw9YNN
2V2szAMj7ePxqF6ICOr1dPi1BhEcVDYEt5X7j2PlH+u3Ei9hY0tAXTEgnOJb3T3M
Y2tGvKstFFjYfCArV8DoFhqJzrZJab+0GWlGecnKjKSpt17dhaeuHXFcRFuN6rmr
4W3JPwR7nMgkxqMit+TQbnugz1YFlBZy154bzzxENR3g9eHZH6FQJ5Y+QM95i2jq
cFjkVpENz4xVf+rfDANh4P3A7nqvHC4ZDvu7yJOVDcayBSAAyc2ztXYS12XfHuYu
EoxeO0oxu4XT2T8Cl6PPxIul0VtLMfEUFZ48j/cleiy4FbBg8IN9CRs/TFinmnbC
8O8F7eXzeU1JzNWL6A1eqIYLiZl/r7qg4gtCtDIGK+nWjA7jcdcoZnEx1fJTS39R
OQtVFWVnJojWmqKHvkk9E+Mj2hODjBYeiRhCIgRPVW+wJVi6OBx1gvppCwhrn1lN
z2wgtN5dSlbYJX1NH/P05+WCRcFIEKiqmUmzxv1NTCqHI51LBLpsQs8YvigxdM7w
OSWB8ADIlENIl8mVl2nU51ezc9Zvyia76DuaiEohrbkTsDJBsKYBTOiP7CXmWr3j
PNifRdqnRwPQS4vqHj2ZlG/kVpY6yo1F09XIdwhZ4DlAslRSY1JOu3rZ9Kf6C5sD
ZV+024fP05uNIpQs/8Yhi8lDQnVV8Eg4lZL3dSXiVlCVoldfsa1kfQgP8mgGBLl0
Z7Rv4EevRNSNvg1MHoFEHeI3lO9tQZ0yt0hKVXWh5fufxwPiH9DHSEkJBFFuW2MV
YVKLF0jLHgDYbmHXQU5XzJ7SBOMAqT8YfRd7/5j1xbXSG+dceMt24NYkwnr303x/
gE5FNmbOAMbP9mvqIPfRtWFr/T11UG+gVjl8/OmlBa5q63A6ECU5EsjgKKY7UKlg
k53+i95eBkJ8YuPT7vNX+qKFVWBtCPhmEnyjVJ7F38/MTpFGvM+DxRMQuTNuwvbu
wCuwcPO38OKsvCvq36G8I+RNYxdOn/Fr5uwPzwlaNY1xflACPMURKSWIO3XxuVqQ
+HAdaRd6C8G29o7PMQ5ASVjHQ8532ur1BNLDKcW4U4nvybPrEOmbYSnZCtf7QwZX
PBNzyKsGehKlfouazznIF2t2VLzhbBKXSgGX1uhUjtFdsrdhyyncFtuWPbDfKt5u
fNowTsNKX/a6HJVWW9FY0qPPtOKK/33WsofEt64Y1lKX1lStNLOTJrwIK4kI2WKR
9kkguJA/wG9i4GYGqimQsKA16hxv29vfbNtjkQ/RrxvSsN9/9XodADRshd5h9yov
ASTCZ45fNjYc9Y8SzJY1LghQIWcJpx3MEcaHUgIpv6x/3J2nZJOGDkkUpacrxmFj
k2rNj63eAyUM4niX/+VaIYEwHKREKCRH4dVQ3c9SndC27Q/0lJ1GysTmukcZ6b0A
DxJpQrreAnEfikLvKlaQZYyn8zw1xiWfyXOdisFEMV7JlVajebv6LD3J5Gyfzbbb
vj5GLvZDzbnFK8fR6ng6EC1MTFNTSIUp6oYusQSgFJkuEC5Gdqh6PjhLwERkLyF4
01mDpbKlsA7WppwW6BgwB3XBpgX6Vkgv/9sI54ks43U2zy5ervposbTYq5VVHGrY
ycJXtSDJ/h/vNKAJy3EKvcalsWvdarqxAYgJBUGm4O14M+GjLgYDF6W7ff07GEXY
tlrqUEyj/UZX+bpPjBpaNDHK0DWai99JV9w/r+dVLH0202Hkc8HQG474yahODEpK
EI8fZs1Cq59vOise06IGdlLlnI1rYjLKsQaD1fkJ8mUIHqv5Jb+mVxgiPkGaffmU
wJC+0IAS3xC9RbXOBPxKg0R2iwCVuLPkKO5EnBZgNatVYVBvjBl++UowsFphoeXI
h6G9IxKInC53gjDKChySWkDLA2tS+lfOaoQWmn2lFZX8rMyvwjLefj3OCcNeVsdI
Zs+8RyWU73cUK+QSjLcU6EdXzUJ5/N9lguGPhgO6N1dSIRCVD8WeH81lCUAOuaNC
ep+40AGi9IeedzISYxzSikZj8T+qz8VwIFaUVJxNCwQP1TLtEzPZLHfo8Pv1Q4RX
NQsX0tbROhZPLp6Bmqo1rgF/IqnZR5ITcSNFroy+HixMtOtPNWNxoOmmdpl4KlGP
0AQysVXfaWks6FWTYUoWgx0cg7P6Zv5wp54GXhq5AyxBVGAOOXaY/vaAlalTooHL
vSNll27mIc9H9Y0qGyRm84U/9BS4fPTpi9/T9vBzHok2RDkEuYy0opDhCwkXs8zT
bpEiu0K3UZ8ZNM5hom7Q8HdJBO0BY/VoJtc3fctrp/cIR4HbTKp0DvBYwilZXOVK
N1+A60wXPJKaAeUupN0l/JLIPkJUa8ItBpqDYoLltkCy+G2qlTNWtxQgX84dcva/
wKBJGzC0rOXyBKehW5rIxIc+c/3ThDOZVFmZJT66gFRrdYFQSgmMi8BljQ/ekzlh
zxpWM5v7QplcMUOasfU1CQYUh0zp0yuuNvreIeQ0yB5h4CzsA0q895RysFco9fCm
N5/I5fqUDcTLgnJOunWGIK2JdGGAyaJR1YAPMXM+szoHXg9M3fjLBvSlRwhRIkXf
F/0IEIA4lmO6rRnKj2vo/4ZHqGQ7wIiwUX9u0bspb8TCUkQRM9FMq5WUBR7ysCji
j2en6xC81788/sdPIV/qTSYzRFZ/fSLEu8ZeSqV0S8ciYgodYlhBZH/4C++WGhxo
PTehtGrGqxNa/pHfAw/hyK56IqW3GmHbJeYwe04Hnz538+2yOWJ6zRmK2n5a3MX6
DC3gExnVrgquIBIk8P1rwwnrPwMb/rD9IzhSSiXSt07mBv9J0KahA0h3+Ddg7HaU
H3t+NTGbJFI+w8B8W3H6DuFQVMbyWC4b47lwHAjzv+NNToWpa7Dntug8U6ktmHv7
3BdE4d8kaZmJwbXAEVvbC57pbvxtShbAKUCZjQLZUzRl2wnprN3fD0pcTXdrAqf4
lTgGUbnSw3iI9YmewnSzY0NwQOSth1GjLv75TMfQ9RWGdceCWVQ0z1Ov7/mjl0rB
hb/vkWyY8gM191d8UcCZLZTOu9+5L6oDCpYTOwltNnzxBRmI++OvXzcoyX3vbc0N
jWWf3DggV14o/9xZg5oSJ5p4mTfI6dFhtdGZ4hoQi4bb8EDqgolb5Ch5Gzoqg6h9
CSmnKGGHOidrm3vXLeBSi+B6CKZYCezZMcp+ZVISJH0b6dgA6B77ciNEGyhTvgwU
Izw/0rv6M99UaKzbCRUP1pVEkaCTYGm72S/dQKHYr9gVhp9T/GXTmEMA3f5pO/I9
fBDDDVZcuodJI63+uHizUQIBjEDr+rfpYcvW0vprsdfrlbDPoGnOnInppyIvBRRv
QNVKgR1O12zj6jgXQVDxQM8Pd7UN6haUFSd6sXhbcvxCX7/1qFCm18UgdvYETYxX
1oQBey82dBOyYKanHjUIBPM715lP6WHPfXoJOw0DE5uLbgAjJDG6PmzzRTMgc/qJ
OlUE9vMUaFa+b4WEzhaNFkbUm5lJreUANf/0s7XMpHGMmr8/bveJhnXva6LZ9nVZ
1W8Vqex74fnoa+5qD2TPWGlLn76cBA5SdcujBGLkAcejIzuqIcvHhLfqlAKggOU4
qf7L6To81whiGTt5SFpsaM0IW/sjWe1kc82dlxvshQpMZJUrJzs6j+ClMTjTUSZk
DI+P14TNoIioFYcBBlwUtRMqGzTbEVc8HKN/Kg3a3QNF9aj/co4O0CiwxvcVAN+3
8trf+YuKJFx2F93oDYl717luMz0hW1bSjGLC70jm43ibr69cEpG9hsGVLEKjDdx0
wOby2DkrmPI8swWhjeT6v4gVebqz8vOMWo1BXjEsBHJRFsOKujBF+2DdjhyhhuSe
0y+BMI1Yiv9DBwNW7+oSDUMeng2/19kGcrkUkpJxQV5q33s4Z7RPKiTQFvgFOc2x
I21WjgM+BrBRGzsp9F1F8IHMZ9AoJjuZ8SaP7Jj2kCXuSAH60Qug6fXw25LTWYlv
laYlehAaxaU6+ZRCA7kfAUdCn79B7gg0CAWi5kXxSiVNNO7+j8MuOmr7tDddVDAp
Dm72LdAam2GpQkUG4n3GeeT6McFuauAbXvFqliFyVirepUxrLhHGvXkKOAbpU3zL
VYLFc1mQqSTPu5+khBVOBEs1vUc6E3i8qgGmcQTWHNeW4JK8Qn8L/KNvc29NbbRe
DpjXwZ1+KZ5j/rgD9j4rTxttk1/8APzMkHtfuiYRCXQ841g5mpy6pkKLbBMk8u37
nJLw5XD2OtRtEWRXMdYHPw4qgc8Vq4WKFtMPGxN+vDV2Jcjwq1dVO8Do/U7tOlXP
hPe28sLgcTDtltFqt5kfG4HWiicS6xCVYlSbC2pZ+4HyTN3CQdiUPj4VP1b17HPK
xvXZ+X2oNkfUy81TkFo+h86rjr4q2BbqpY2Nk1TjOVYQDxUcZ4wB7oNS30MlMLWA
uGmBocG5oxWFMulWYT9YnbTf1WOOividtAeXm9xTJX+lfZKVf2i8g0poAuOmCvYM
rHB69s1WD+6fX9kv4TI3p4HanCz2pGA//ibAgsgefHyUh48Hur4gh495oms4h7LB
TsmzEvz666B2FA9IwKRHVPpYFpROSXLJF4gmi87AiZao2snpNxeGMHh/ah3J/qwv
eO3BCqlHgLFBaxCqT4AC2V9RhdDWErN4cl0mP3z4ZFJjHDVqKHW+QVNcHVwsQBtB
NX+x+gOqSBakd77sqqVcdp1rIUMCPLvKuViB+ChyhrrY0bZBK+lFcucPU1uvTtPB
3C0AxCvMHoUb8CYN++5qGAwkHl+DEWFxooghp+PTb6oIFLFfJl9EIgCkXVHFzt1y
cStLA8rOhV3r1mIBuGYhdZk2ZXY/fuOCSWUNUET5qUsaTrAmPsq8/uzZh0r+qxLL
4A/4j0uI+acISvJN2ZDf9SlhN+h/8S/RbXQBelEVkloIMnYu/eYfmVKbtO4+BupG
7IXtZPJECrvrUpR/KY5jjRqN5a36tcWW05BRkLTNDAXTsf2qj8UVtJO5FU7DmiWv
imYtdn3sWNbEBHWgBGxsM5VEJgcA3zWjWKY2+uy9w5rlBgl4C1PnSwLXcqckFcZZ
TBUotu/m69dljpvzBp/yWV8h/zPIKXyrE7lReULd9sLMcnlCtUiP2FT8fqTb/tQL
wI5NJnzJlIrtmongnY5mYpuMXlsd5nsu9NZOHZa7UbW2xmRCcLUsvmM+UBBaONVV
q67rDrDx1Yiu6RNxZX3SSl5vCsKTC9AiO6eX6pjgzYHY8iobHGe6fAmdeRXLkTvy
iZGFHXkhqi9LvHUm+TIGjOlDh88LP3L//7HDVq6H88mmeXLOeMvBJq6PZyqGNxoZ
K3LvS2aigmS3PcO05gi0Z8gwjr8BrcrIvqtBLXD4p2psUKsUW4tdMhavcyairItR
5ZC1vkr7Mx7ufPBVRvQ4mAYbTgRmpRrzM7pvIUge9n5uxjLwO5E3MrVqweQ7IDep
2jSxXRLILTi8PagUMVEsrNCzcB9oSSEwt3uXHYDo6Hlx/hLpAUzq9r2i7P3D0rkc
XJ+F3Zd2nL9oJRLUzlqnUlALpqI4qZ9HdHXdZBS0ZNWbaBLMfwDInGj2bXcyB9SY
Le2Ho20Ec+dMj+OYdSO9Wm/rACQblGuS4uHyouHyGoKy7+StKltRiEZLReKaxZ+j
VP42Gl8eU2gaEDpuIa2Aq87tN7vMvhNIsRANYqjlWUhjgnfUr6+Ia6FWhTp00ZWu
tA7pjwaJX29SeJmEFIrZ/c//edCKSHvaPKq4yJy7yq6sYTWmzQng/6O9ni0pbmQe
7qqvNCnYc7OmtWdlYfAfup2axDXMoRiKWH8XTK1dEctK1ZT10EmeK53i3oJn4t5G
ARtSLubId7jzQbRK4lWYazosrYpFK5v3I8Lh4Ccc51eHFfZKTn1wocSOJkOBYDda
ji9DGoMdvECeZTYqLFrL2Buwdvg+z/FlbuqWWErBXBNFWdCdFak+Yc5c3rhp6YCm
iYUMKaZs3JwK110HKqYjAKurUAxQsrefdrjtYvOxkUwmvIyUaIhaymoLnaCmFQL4
PPe+awNKlVeOZqYKAi6KhFihD+N/55YG/OBg1iy5mZCW/BDczff6Y2spQbmwLkIl
8rFPZDrL2rxRniMBV05CDZMu83O1LL6hBT1A55VdTOJtMsHJkjaj21HNHGNxMQ1a
emXZlBjdBc0/FRAvFXenvoMK6Hu3+kTAdEvLeHrIu5t5anrq5yGBEfg+9BG64F+R
NafujajIIHc7R9FRPEA8/pNOdMmDlbFqYXM6S+y+YyilbE4xYxD7Igwt1c5KULMr
3wK1vEnc1z28zdyTqbztREpRUIiDNI8j9gBSuQ1yeb1FMniOR8aKyiby/j+ZaXG1
AWitOzfymNSTzfxXW95hydjgJMR5pQAqWNT/fp19Dwbf7iPXQnXLM6SUmTQpA4+V
ideSBi+ka9T5KeEvfn+IhhPMPMO7Zn5Xbu9TxC6DyopQYZ2JRsR9pYWs12AtJ2V9
wd+P6hoSfkAJW5MgAEZD5qyXZpal217b+V+WU2EkEVsrGK9AMZKaTzMyxILId2Kp
aaHN65cFIUb4k5cQ6v+zZXYc5A7CMDLneQhwFXtjJMp9aUWdUVUgyFXoy4ZUZB1g
qPD3sKjDdGboskGtV+SLyIm1uKhh5DYdGSLQV39NHrB4HkjNE5/OojWdHVLcSh6J
0RLp+z3zzEIugbibhWbuMNNdbSDGfKikuXL6V9aQBPJ/7oUbaONxMlF1cd3+61Yl
gqaxwPUEpSqmhW+wpPFgUY9eORamVstaZfMpzrZ7G7SLJkHREfkHnggtv66M/82O
qxoObfOgSExq6LaTeCV7PFz2GPyHS3xgmGNgwEx5scleCRkVrRHGVx732Jau3nVH
PNRZr/0h8XjWxbcTjuer+Locg32HXuLS6ThRcn0J5TVu5QWLph0lM4rOjwcRjwy4
I3BhwU6YK9yUsBmKmbPZuUcRvRuypWFpDP0jeH0SwRby2lN94DLurO92AqgoYgXU
dCMjM1SlOgDAHk+8pgW5VhcZ01K9n4V1VumqtSsqyvioVjZO1RR6lOJJlcJz3y+T
ndweEUmPtBHKWeEEbAZrFKWoqkL8kKPQ8Ym6/8usZhYlbYbiV1Wbnogj0nAluiFG
dnzQEDG3qZE365fduISkTSJdzZkK8tTS+MHAhbEf56FVsvbzmGu8ADMRnbtg000U
dnJ+gU837BYsZhWrTCwzxI+c1wA8+im+yusI9dMVjJNt4Wx4VYyarBfHpyuF5wm5
kLhMFObobZFs42yHppc9Qe+Msx/wM/VdRau8fBn8wS3l9iF3WVTD11Pwbh08/261
6RQAbyDagC3pAyvW0CVAeOmWy00109nO1oIMUP1gkw+yo0jU7ua2xg0iZILK1Xml
FjTGJjbjPYZtS+32+qK79GwCmKEW+7wMT+aj18CqBIXhfvmIW2kPG9COzN2CbaUF
JQqTsz0PgxQPowuFN3DzJfGg3aCqawRVBO3oSUZxW5RsfUz5GCMGjpCdyTA4Ludk
h1z9p1zeai5E2AIDnPEEuYgosPv/UpVW7eEu+io0VbNoLjWXy6yZ7aQNVDVwDxru
1qfVUpsRlI8aRbQrQ98WAw3BzZ2pSn1ivH637V4iMnnVh7tsCDlZDwHvONIPF6G5
Vvf7rF3+Xs/ucIWGCtRVooyegDJWXQoW5V+UZeVV9ouzEoTHPVNUncRMjrr3kosP
ME7bC1SNuARdw6blV0xYuv1s3rNUZ12ataE2gz290pCH3cyhsHNOnR94LKWxo2yy
Q9V2VSJwcmayK3BT4utS6j/0xNZnZICbg+YJK4FBzkAeGA91hG35r8lFj7K7lo9l
9joF4Fq9R2BUPQXNKSiW/xdWRLj9+oFL459UGxJKjSvaTUM4aStUdawqkGiQbGLm
5Uoz1fBXq1Se1/9rD+l718qLCZHeRl4CwF5p/tc18BO6egHo1809RkCiUQ6tsTA3
UIOqAbMxydDv0qTMvoZxaJGJVqdDx6MzKHJOIJ8qvtNOpCae8il/tgs70qpPYSdL
MCrv1606aa1y+xN+EvZ7mjcv4XnXEuVlKuANlVBqoBuCgQC7LhGPxhyO8oKaxHW2
dhbrWC7QI1ROmFE19Beu28oJktw54zq3zckphCvxqt3dD+VUsX+npd4AZoFSvFV6
L3MlgBLUAvukwrDqaq5GaNKhBtKHn/s7EI9Rr5esAab4XhqCOKm9Wp/ERcX+yJo/
eYGvpAM5lQlGmwE1ujJyWl3x9bMVR/09Prc1vIhtcwurRiv8ZhqeRC41jqgfEXFV
GVFW+tSas1YHlyn1+e/GGwW0biyi16hXMv3Gq6kKcyS5i4lEeVEALj0cXro5LoSD
3DLlhDZr89u3UGRKqxnpFvIPi40toXs5K+AL2rvZpcSS+CvXhLC5eYL8pLvskLbC
DLKNSWTwrTvLfQMoMnnt0Jc3q0TPhi3yxwCRfighBSgTkklo0T0AbdftygbD+lwo
DxHBrsJXBaWq7kavazVo4rwyWdtM1jBXA/PTctx25Z3c8pJ8jZ7dF/UqKChy8HNZ
yG9jID7GexPSjVmE+57d7eANGdyQtLv4jk5fHT9BO2iq33/AIvrgz7f6NgAi0iGI
VN+9nqiIu6zCyQyfWQ5VTgJWbGIf1Wq6GOjIIMkMcoa21KLiA5vehLW4tAASOgs8
siRJzXDLXin+DMa8M9cTdB0kKSHEPZ+mFAAV+pDKEqy8Kp2XQnw6Qx66LYvPJFwt
dzF6k9FJjjiGm9F3g3XNmsxq3uXRZhEO9PcXTnJa6pXvbfHI1C97u4fe5SSjdplH
5P/y6cl+OwEpWK25weyqtY2CDr6EZKJtQd7QZcao/nyZXVJA25R8zGHcfRU1NZC6
sk27B2HEY9D3RbV+vFRDYfdLQ+L1tQVUc/lPq2gC6Q1GKJr9e0bk4uLpwtZK4/+v
ouSAE7fiDd01FD+/x6tfh92qRGVdIKswB1TgWAhIMdKTgSiP3H9H8/9gycCPI7Uv
pWGD2fNOk2AGGWqo6X6JZQhh+uisxVmPi+WBF+JlRTW4IXN2VC1gLV8xGuPDdx6C
SaT0tuKs+RpL2zJvQr9WUkpAwCegSohBXKgfZvO4SOG/DZvmD9WimH7606sqb7Rr
r9fcf8OIgr3Novuho3UANmAGUzXQ1+FFTn9BLrRRfVYqiJsFab/b+mPGH8u0MafL
tdrPka+uR52/C32qZ1hWbOnBVytyS/pLJjvOWtSWtw1cnNc4HfOH/cKS5Vy3YXK/
CbXBDb4NmZ48UxyKNsCySgvaQMQATRlBkpq85HsDf3GGpLk+SLTSD7kgYqF81UvG
slZftXLG4wpL55RenKU4Erp7t39kH+rbOSTBAsUQ5uKT6oIjLFnJISaiYYDcNVjJ
jLBKXxdfVAxMAJ24kmpYXVUjjW/Rl6uSS2dU7w6TSEbMCBvhiEJokvuwcTttbveW
YYg0Rx8OzOy373vN7YfHfh1Zo2+4RoZDe1EqSxFo9v7ZjAAF5Vg0a3J/rHLqbl4T
b5LBLzMz5w0xNp5G5g5rp0onkKKvKIU/RY1zbJEtvsthEbpNgBKPYy9Lel2Zq9tu
LSYirtIcJPVyFbH3Pna+l2/uwvt44mmCAI0xCIWiDCgC70g8CFzdAeTiUFRxJkmZ
bBNfxREhXCf+h/VSxoLuNcWy/GOE5E/qDCXIIW/De5faIK4XaaMdVbuXbKe9YXXT
HDLpHa+lvUHKL8xyZ4C/NtzOs92v0ifqv5N6pwX9pjTIOQpQ1i/eATpZ26Q5AAId
J6hzKivQwAJoA4sYyrp2JXG4SW65RTXdFlWN/Zv/qaMGb7eAuefcEZd0QHa5ooNU
iP5GDpgNBdWR9qSqQYddMRipZe051N1LRxyJHrw5sxHM0tEoIg/AxSFPR++40hNi
8URhOC7nyyN6tcu7gRRRPIwsNI7pDuu+qxrfEtmRtVxKzgAbKQ8U0yWMFAjvs4Er
Kc5Ex8cgj4nwxM4F3+TAn0BOZWAGQHjwhx26aYTA7HxewghxIXDU6poTY984+FXp
MF75airFYk4w+0NUe/X+hzUakUO3yO/6XuQaJ54VLTMgPEayFjlcdyRM3NKd2TX9
hoVK+DncpQL+iekrd6to/KCi5a6DlNfOHWnggQl+LFurHpNcomr9hX56CHg0PDYf
t2Ucue97AdPP1Ic0C6jVfDFEYuOtIIINT6oxi8kagSN0mXiEtByh8NmTKMyjxyvz
pDhAVGU1PDcqNbhtMeVrp3InA+XNPGNmru/0GVjFdpRXa+pV508W5kjjwJbmEZm8
V3KHaLXbIH1AtTTSB9qB12aDugoV2M/0+5/6wDYu6r40QYwfQz6UUgjIFDJQpRyy
jofXnae7dYF1fDW/c9XCuhb/PGiCwhStOvsiijE14+Cb8UJ1XsGfuU0NFlgLIZi8
G3TuwdyaxuWzWmDeVnAsiRSd8TbAhIus91q3auiG/3uGctKDYp87bmLwPP2Js8bO
APzEV5btTd7WXw8eznho9t0UOZuWSjA0eRnBLFW4akdFRpxgZC6ghqCwhI4sno65
lY29FamlVyJL3+jUBxrMghj2Vow15uxiS38cSo6Xl9N9HTrLec5ez3O9zFbyxcoX
rtduMJ/AwcUmCdXYVk34W93rBIVBqT3ajqDYxBFyrzQK2XC4ypQykRZC/i+MvzLr
7Ic09qSzdim/lA8XkC5U+wlCU2tQAOo2bCV6HGTSI/ijgiguBu2203kF+2txpaXp
R36f4Bfbuz2LFyZzvwxoHQEAz21JzliAssmHj7LptA2Xx3oYqWjm+FcmcSYnfg2M
tpvAFcYdvI+kh98dfinnUJe0/5JHk5M0JBFLeFXUq9CoeP0tf4qX3sU3tiFOOWzW
hL0Hf7ayqXVxponULtxVHd+3ycNCebJXsYtKvxXAaIkiSbkgDDzClnEnToIWYiwW
WZCf4BLwnOUJHuTdKndo0oqAHvoQ0ryjy7BeRYBIp/ZR30UVq4wHVR4cPybYv5dJ
dpGYYtTIBCR9I+0Q8cAjwjOBEi4jgwDOM0If72UGw8oOUiqLNpekCvgMIEsWoY2V
DQ2aaVfAdAxVLZuELXP1nRd+Jt+6cP1m2jDe+k4YrNvnn1a5y4tf3lGeKQqplZdG
Ey1JUE6ZLOydYYCnwC+PE8pfOGFKTx430Graq2roS78o93hTueCgTBfY9+YcmxTb
rx5lCQJd71gNtNrcdAtuWBFdcxs1AnfDe1wD0kx5a9+GUoHGlJcpsLkLsDpZKzNz
z0jcOE9mxOsKXTdArckrZTs/NKZpDKFMIFCRTUuKKNehffz8sCXPlxC+4/ceKM7k
D/eyoHXQh1gMMPiYqhyIqm72Q/PdUViE3VhbYbzjf1NHP6xE180tpTg1iqqGsKxM
a1S3SwoTyYj1aAjD58jXyXhaql+vlTqhyYTZoGdQ+QOm1LkiU/d/AzuaW3EAPL+C
RS1EHqjJq7ir5jbjvgImvDRrnz5vESYxvdY3POYao3BpqFVpX19PSRNQEBwTu80L
CLqTbVhDP6eQMDypaykxTXbgQ+u0Wy/Yol8MU03ojkNMOmhMUhRqb8yo4hYV1tLp
oZNol0TzZJgNrajz99MLL+UtowMV0HHc5NiXADYOZYvxbzD+jiWdRhEdISsgZ6QB
Bx4EACsONfY7D+KGWEQp+ZjRgfnQfEtxYmDphh5IKfrZEn6BaYPyJX2w1nZLdgpC
iSfNoiyNXK524LQThnIR0cvFAX9aQGRkce1HJJlwETxStfV+nhS4Znrt+r8XFQy2
2x1tYdimtL2xcdQn1dbR4sDysSMX2FqqeABtpehZUX14IM37j1LjVdy/HfNhosUa
K7YrRFzatgtL9xue92G2Whf2j5qcNMkBS7Zp9hfIN3l7UKStJGv9P/e6bK3If4bh
XIPjkEKkxtoRRns5AAs7bZKV56we7QYqC67Q+oqA15TA7zGs0848R6izOEaNTjWb
HDAUQ+l0OguPt7qoo1Yo3sM/qgJducm1f9lFreiNe82BMRzfgZm1LnnhBqvP/SAR
Q62Pe0b5b7VZJbwTi+Y2EN8fb8ARZyhNQUgHoSsTXnYmxvk8yL3sVAO71l39fY82
Fq8ydFaz45UzhPlTaKHSQht7jCEJEfAEUZpJwY4mrYESOOjchIMjSd4vRuNCq3qh
QfNM15GJcFNbbOk1IR/dazl3g0ZqbLtvDd4AGooAg++5L+QLrCgGVswqgCtl31CA
of/pWRH766oglZL942xVgVuyJPaFAfKEp3/8WwmcnOzXavrbvFIdhA4p3tnIznWS
KvWEHiCrQ0iyZmjxTCMoZR48em3KNX5hM7Zxt4KSTr2jNA7Jo6j2HSgBo0sWGSwj
cqfD198dvmpclg6xto2I5eRWXuZzDt3XR9k5EA4a4Xm+L4Bls3+DyqM2s9FCfwbu
08JnS3jcsf3iGsgJZQJH4wHSI3LbY+ieto2ai+O/LHaBNlrPR2lxUzX3Nfojho1n
KFFYblvcv1f1hMqBoKiMAT9eeWksgZw7+cG7PcGQuGJTyeIu9u1kIjm9hM/lpM9T
pg4HVVpdvLe7D+5qsRfIzV7rn8O/K+5eEOk44cllLef+E+nvXNl0YBiYFpZyoAOG
uS5DW8al/tPl2FfJJpG3PuRUblDy6GgD4nyhom/gOXIwOcQOBHNy8G+gmoRI/dHL
K5pgCJ5jc4xvcJGzxI1blaN5y1/rqzc8mB6wF882bhFRfWvXaZyGV2rOwg8DEMMC
HZfaFAv5sy+uHwN9DthbCwy0l2zaav7r1HDJc4uDJ2ttowumuKDtXWXwhRWns7Nw
nB2aC1liWM+mGt/qzd5JnRRCOPOKiXcAp0UebYWP5C7+42xmWiQzvv/cnjlRX/un
XPIvQxnuuW46dVUmrL7FoiRJQnqw5Wz4A2Wi171xcWZB9VVxbkWC551qdpnyJpxD
aNJNKtmnNGw1ucAI2mBTHS8shHhc0lFwTmyCxMC4u2Qzom0mEu7Z0vSFlJLFfmS/
9KVCbZSmWnOWcUvPp/Qgq5pSnhTKLzwcJPomIn/FOJlq9liYU0WX+3fNnIqPWKHT
UrZv+ZFYK1OaQYDCDm6lUq9DE5HFjzZvtMHhi9mvspFVN6RkDs7o8kd0VkA09T4F
KBwOF9Iu9GhKtgDuNhZirnNnkuGC/W99TBVGyKfY57Ven8nyCR05HlqkLFOl+JaT
5acGXQIhVCPWvsgKUVuf8vQ6qsQJxMUdwijbKTFEYcyvWliJr930ZHs2veL1EDIA
Yl19eq7Yvp1NrlTZpm+CruK+lhSboyVcqDCeo4pbTB+99X2l0O6CcQ0SuVHSN28c
B/Cgg7dfFheZYSPVepmzXQX0loc1gkP9ROxR7qn5GfWE5Chhp/AECBvZLjjzYruk
7JhgX+xRD8RZAIshn84fZ89Jtz4qjeVm6C33l4VDxI2rPUH6TH3eWGzXUzAuqw2p
Qr4YPjrK7K2BdXXwM1EDfpAMRcrnQOzLG7x0Oj4Tg8cbzV6MB/45KJWI9xqUmC9a
q1FXTWsVq6DPqdzEMMigzvdhtyg+ZNJmITEhOcuTBb4iXOBuoiXn37Xl6VxnahUd
bxiP9jtYgEST3Jz4QCigx8w2EcFPJPhnAGae2+44swuwPPhA90e9sLXD0hoA2+33
tvcTdj+je9F7OfvBvyC05zbd14MAbdKBMz8hO4Ppo/yMJvkg6BHRn/nL4gR3yFDb
U3SgCbJ0tvTPxRgEnosGBka58XZEFNgSED/DIKIrvlkQ0bF1AwvD1/x/9qh9iqMK
Vr/548Modz/1wyMhEE1el7YAn3x57tw5ykIzSYeZ4fWKXKs08MMwm6zXd9GQ4slW
DJYGRdeO0/OuNdr+ko9HTMj8Z0BsVfcBBxiS9bkb+0sF7TBRONNCTxWTbrBOMHEn
AV2oV1EfIOg4MdN76PowR6tiYLVfApmleMv3KttBqLoYUFd3ug21FHBdkKf8llUE
/hgGOfjmxLIodcmkejQTXXlVl69AJHzO7B86MZVVMCINN58J4KkzwlGbTPc0qIxX
KawH1LonVS5ccaO67LyO4TXKpWiE7v9UhmLUWTArtSLc5yOlEH/MqwZMOYWkMKVa
rbpyb7HT+W2kgEoBEo9KKt+rvSSM0o94tR2JBeNEZ/v0YApwJI9LMSGSQR0Sui8E
gKQZCgtnZxvgIKjaih8y77hCN1agNVJf7LfzBcITVPxnoMfryu1noJaXNYGTi491
Zf9noqwNi8aF0z1N31TvfjMSNVoQIvQxdfHFKv2bzIW0e2X11JI7L/yxr5SbJ02k
/zWpb/fIvmrd33aDmCwwA/5LbVyG5ykU6hdOSzru0Ff70Mbcc6QyPxsi0T6r+JfH
HKG+rhCkFX+b6pCWYjR6Icwb1lnTbALmAo7H8NgqyqpIeoyc5zVupX1nbC3Ic/QL
7AnrwH+PXsYCVJiH6wJwaEzflbyU4Irt6J2eFNsDGQEb67+k9fmLg1UjQv+Yp4a2
irX8GaLpSNWPmpbolS3E0Yk++aejqqN/mYqUAWL4RZyGJcYlOCH2MXyoMm+RTLcb
j8GQrgd34pNPsXS8ptJ9YItgqFzd/M4nTEX0Ig7FL1mxKdIT2rOBI9FuMTig3eBJ
Emj8o2qWc8eGfhLqauKi3R3WfOwd4RSmSL4hLTs8GaMp5DKVLWW8VpdDSaRvel+/
xAY9paiLNdpSkX3CIN3VXv/tUss5NRUF8lWiHhy8bEX96QIdsLg5HKQuXYAXxbLC
ScDnOdg/53Sj5ViySEHf/2wuMzfsozOF1O2n2XpVmcEgRA8RbEPOKBxDOdODEUlP
fFGdZwNZAJFlI5AD5V/zCCJKmNUD4G48KolboDAUVxGJ2GYABiqYoy6EGM9Zi+lp
Gcwi01ex5Q4xHqD+u5aC3jqqGPzXDsiIalPhN7RE6O9JxJkXRUubUQSmEuMdV40e
DB3/2/ucgzE3F1iB8p5c3m2wlJiL4HShDoWCQltFEwiBjLPTQJgFvAcaz/yKKFdX
5x6kcwaHoXrHX5co7O7DW9CjQ6n6lHQW+BtbZlFzShrHtbsbVZwOaZF6DPUYSYQ0
Nm3wCHClBV7tLxdr5YYFWbOyx0g1bYEDNV188YN6pcrU3Jsn+v67+eULuQQDgj7L
dV9VFed/KGSx2YelIqrnC7KvHRrtUFFp6+QYri1YCDknjUwCc/We1GG0xGHD5i9Q
gIAoxdKEahNeczwVOzHzfcD1Kqr+XNMtY6X90uRmpD93bOgNwwziBjuvjRycdoQT
tbgQZ3TuUtGdA8H8IFn4d4C37enwzswimopdqfzXQDHbQ+BHD8sKvUOF7UHuzeJv
CxllgpRAv0AnedMnQhi2BMaZnT2mNlJWNbSktCXIKAOuBWJ/6HBFxD4BkdpYAqrs
6Q2o/B+RfspLAXA11mL9iDzg+1jRY+2oVUEiBwDoOvd9LkKjZjLNP5Pf3x8SN6jC
Mn6nAHPdg14dd5lKak8osgCdd2NeZMBjO3+915+DYy/VfS7lh2mRSZOwIWCL81dU
h2UzPsjLIR1fTVwndOalKYfl9RSF/+JtSrxwB3pHZ3ut2xE2FOyAApNN+pQyxzsp
RjW8uutlaJtc7pl+kuLWdZoDYa2ReWPst0RsXR86Me1QgbdtV8CfI9xfTeMzJ/xg
12o3XGgQFZD52jOK6gPfbVmkcE4yiyPJ4RafM9oQAgG50bgyRxdvMvt6NhDvCdCn
YwynKGDq4uPul1rRYDxML3cXavsF3gHwcB9V/rA9DXH9uUFgBdskDfflCuebWUce
wj+q+OHp33cMyGFMsk6TVaMbj852J/igWVTiRN4no8EG3w8Sg18QdbLwefcInXcq
308rI++xMd+wqNlGWgGAnzIDNHXWnQJsKAxHY8eNIFFkYp4eTtLgX0W+z95LDfZR
/bhR+npznziKg1kx+2UFEVm/8T/Qu53kOz0WlrfE8BNF/zXoUKnJUpFLJcH/a9aM
NK8c8SZSM1lqLOwSRw1PiJEryOzilY1E6fCgxiefxvw3w5ADsZewAMklBgz1HDFb
AwXnoryTggsfwgaRQAEyCnnqXBVSlwJwn62PqoyQSIYAxtqFKVJW+KktCxVv4f8t
VSqrrjiuiIpUSsREEIlpCYC4f0k8zQZwjB0sQEhJJ5+CjUPDm3BS68D6ES2j5OPM
0epIx6BswupR45g9kRABPD807TPSVZ+sTx2Y1pvPu2aJoVtwJQKzMbtGAr3W3xHa
JUMhDldnrYzaYCeL+bTdjcyIoaM1qlA1pWSvmzSMkjnjTawzGwB3rkJ+zEVZrukP
F+HE9hzbMmEZAF5ADAhrbz82ff2VO6g93GybXlpR1sJ+UvRV02wcSVTXRV+kG4Co
ddHDcEMLiDq6bmls8pOmQDgVBIvWJ7ago8rua1Foix1zUVVlcBu2N82L+P/PzFWe
kOUD2CuIgJkzGxDsZbJz9HGxKtYUmb4WedafzvRd1aXpZIAcZzkDW1AfvDSA/cvs
OPRoTmDK7inL6ri562Zu/iW9jD8KWIbliOSnqdHqmXyz4LZs5OUYbEtEfgjm/0Vo
KhhZZPXz58J3HKBcc9qNchwRAWxNujz9YLPUgzcraq1Z65GfN39FcxxkiR3JNR5P
hCg/TCJ7tcTxftwPoVW/TpBI9+WogmbJ1A6FSV4ixdwd/+JzqPCQN4fgymhYnuP9
fv0NMjBCZJYBPFXQwuo3anO0rLN19uTDi+B0uCPucS5W3V3U2QUv1CwQrOdINfNs
goaC08jK+Qw8pdDZ6ySdnKIcJAgsPqPWwnGG55Gl47xUWNz9M9qaxmMjBt6fXHWm
3l1LaIn7jKtUdS98I3HmVSoBy4rw8wh993Wg9lOJgozXH2h+Amp8kg8XDABY7LOA
mns18HfYhJ+12hhNPNoqf+70zUESzyAbO6RGTa2sbEkfh+Jm1R02rScvONU0cH8c
afzEHEU+uAUsl9826y2oCHAKy69gBMqZciS/GR0ajJe/rWnk4l76B/yHMAkEJ9O2
7KiVjtCSE7bLP2X1oKPvleKmK26stNYixcu6SAE+iWdVh6mtZi95pZJ+yNYByznk
Q89eJa6vMagd/o4oyCmTFpPvuX/FrTeGI4SrfsolAig/Jf+Yjh94+KlPRW5eu0Xo
fosusOh/TqUaNIvqbAnrQpoz/yN86NxrtYBFv9fxOpJfdyxjeNK9RrtjSGRiPIBN
acuU3uk8kJvkAoieHsev8zk7InMJ5tUol8VvtEl1Gsz9ACr45dCbMEDW+K0hVeB7
ewsMBuOCkDi2pheWqKlxQzy7w3kyW34LOLrBdfv5nzGPArrKyrMrw+X+CsmQGRp5
ICQuYHOncQcVXDfcNhUB4KE509HsBDNm+JhgrnO8s3xba3MofzvtgJZtCKzRgTKt
DgsLUhO3VkoNdeRyJyEZC2dB5OmFUXhpBZm+nRl5674H/vV9n1GtwxlrxswVxzYB
DNneo6OE97eosYNEXevP3RNgX6BXE7X8rb1Aejv41CXDRgXPuAH5EVsnCb2/3tgK
S0Q5JAZb33CMtzHDJWcvL47NqzKfZfdE6TwwvTMWrg2oVHz8K1t0ry+g2dxi/KVJ
Hyx5Oa1hxRyfQvTwolOv8RTuSHiJtvGPeuiochMcPXpCa/OnoiAzurcwbrJeR9J+
afOvWqZLuLxvgQcg+iRPfXPShYfNmhZmrs5MVrVHPcpfoQXnzRKMZIFh4r5lJhng
VrE0ulqsslY3icYKyGpayAfknQqKWNcO4GbEwELGBS5TyZWilwHfLGOJjkGxYJqO
4Ill1VowGx+x/m72XebjB22YIzmx5b5N0DDpCklMoMYLzWKCl9DT0vQfvmPToUa4
+XfTST9GS09ajglB1uPGYT0lg++ZUt0WwZ6mX9XgfO77iBOlXlCBGlO2nt51+uhr
iMqJMuoNrIEyAhB30evdbSkW0z1jRwa3164kJMxj74j0nXGhEe2N92cnElHXpsHy
5vdOP2WAHXZ9LotnV9hWtUn4F+2Ih8HmByz23cAkNqmnKOUzxv2uaaq4FjYhA3ml
Y9obM+TJcb/eDm1Xgu47QcrYxPCBsbPyZWRJvJeHtfAw+7OxRYesfZgYLaR5i+fo
XYbkS/uqJy7wevSai13In8ZmpoWO4h4FH/TkjgCBvhTL1zLfNuIj0FzgYwVBzktM
AIbhb9ovXaMXpd1fPxlAysjo5CwFrtExqXb12r404BYfmjlYoUUPurWPm7AElv+g
SDZYtJHHFhaonJlxHMTl0+olyfVTHKtCzAccPNnn024rn06eiS2nuFr6otJ140M9
kpu+7rhuNVZMCt2pxXYOGsNNnQGkxK64+G+jULBFJ6D2OG1eiXpACx5VLc2JGthU
RS0mpDFt/99wAnKar3X0LSRAE/2IK39s5RptPUyLmGmPywxtEDrOYht9Qr4vZUx6
gVO/PZcFb99kQwMate76euIsKmAYZZ7KPeqQhvymT8z+szMfze86icTBnPmglef1
ulr1C5K+oDx612OyWS+N0MESkQkBmW4VVMhDgDL22or5ezqevb3c3uGsl0IHBa77
mqURwf0BzuNvN/2iOX5ck9XCuC9gBw5Z7DRqeppF/OT60AokeY1m54e+fUdeRA8i
vnT0Kvhx5bmnDzY2FqCZdwWN6PdR45+sURiAjEidBqcOIIsptKtsyYpj0TB1Zsa7
ozjTNSDpKGugxZrM15enoLyfXn7QJV3GG8GIGzAgKh/138GULnyDG/DB/l56gT3i
9fWVU5utyk11TMXb3V+X6fZ/t2gBMHq5wCfo4xCz/69sZDeDT2wwmhCz2pGOjSuN
5AZiCj6ox/ss1AsRRLPYNzXZfacjjA1jMLaZwoS98/nsPhLcw2UM2kLRZDzAEkpt
O6dQVVwj2Gzfk352fAzSMVNTcW+eYvDtTVNxQgcI52WcXCqsppGiGO8EyTeVRbfp
lNvbbE+HjOpoiahbM8FV99vxj4gp2Ugm8KB2hJfq8Weww3sMqXdsUAp0SrNKfiJ2
klzef7+6uXzG2kxRelwhAuU8EFhJ0bZDtFeSyVrufSizIXMsbqOf3esYEvArkZ7R
G68A+P8RpvSqDcniTqoaGjrFh0eByQacgxXfhvY4sf+y2UyI4lOshHlSdBJZg0kO
Af9ihtngfmjzP7AwxJwGkTLJPErJWqVVzZ9Pwy4vJqilhdZXxij7K604MvqwKS61
nJ+aRmYS504dMxOUFhQteUpJBsQ36f1juGG1klqVgv5OTcIizDS6N4kc60PJ8oJA
OQaUoLOy2scrvo5GP5oFnZ7YpdziEgYQbrlGWbiVEHHbQaatXZmM5cT5Tvxpx113
6JSBo4DzQ4U+GN4eYwircj4FaSrp8+EWy1soSK/vy7x0UFNa3lZJ1txnFN0eQVF0
QI9hr+EOjbqrcYCbMoYCpNP4aTARm4EEg8iHQQ0NdH25nQ7MUPK4giYSxQUJDbw4
NAySJUnPBuszBTuiEEJRGngUZjOviFALO8pot/vcjn4+cqmYIQ33tLQTy6u/y+MZ
ByQdrzjP8GiQcpd55FNrx7u6QP9fcEfHTx19u2Klqren0nvDOvP5DyEdAsRFhOow
Lc4Pl4MDQVYRzbtVjfBQZ7eZYlxN/MDvcgUeWV5PQ407uubhGK6icdlEZO6+6sfD
cTWILTD2UkS/nZya61oEp2iAfzdmOscwzJks2dZgGWEGXViy9a5wbbD+fW1un6wQ
2j26pWKFF4AirFsjFCPb6xfsNxvS4YmS2YqwQIzHsots6Hmb1A8UcZt8DRjOO8YU
teTXhVxx752qf9JZby/O6mlkefjC3bmv5sW/26lHSEk7H1DW/hQvhBqptGeIDQPd
CHNMFlkgBrh7zt1EEnARphkAbA5qqXkD9KHslu7yjQdYo6jikVCpmeDMsiF5R3/f
npe9NKc2tj5XEr2sW3J2VLnCnYJmL7VGUGxjRvU/bALl/BRvW8tXE6z3KbDg5WHR
zm2gNOIBIIkfQh+JIk8cMPEq+SfXCPgkPKVmLKbxDNNzM9vlaeEH9GMZV9CkG3Ch
nKR1eS4sa7wVBPgrc89ieeTWa+QgsqZ/sneOWoJeYBGUeLhdl2RxAh2YO4yl3vJM
t9xOLXWyb9LSb9tmy6+W2z2dOgx3r1psGWa+Tm39Jj9ML+7+L+jI5f6HV2vS47yk
b3ct/kUK2oBxJgfxmuOy8nqqI35uOommIzIXvCJMs12K5+lTjew+snvRvn6w5yHP
qjIoYSsra9vw907ozeSYWM3Z2svXwHG8ChpvK2FGXGkbVJUCOl5TBQhZ7NzOYEx5
HnIToUS9lwA9RHIr6JI1ggMgrrfZNy82Pgagwj0uj3ZqZ81Tstv41QTKvQ3YnZuX
bymIJhqkXaXG2wad+E6mfw5uou3UWpZ7rSo1bsjJzE23hJxb+e5r2ddqX6teq0Je
FPZsiJGgBteairrXYCryDaJAjh/U+icnXpMkAScluUteJssaYxh43Xhix/fIeNPc
PWW4pd4cVTkU3sFRBkDEehtSZ9kZFdiNjneVfHhcpVMzMSdsUT9MlqEycRV25cEE
Qf4Og7KKC7FNX2ar0ddnSzR8kinUrZmqDwc3t7Xeb9uQLd5A4Id12EB5Y5/TzLr/
7VkbVL7CXMG1omc9+Tf/Lt+sU1Zy8DPzBgSHRus+dgUCqyFk8CNHUB7kQQbwHTwV
A9ptcJN/hQcsriHUz22+NwfdXqBd8Ywf0QxO7ZT8jLmVCe6PZxoFSFBOcoiX2JY1
n4VVxWoaYaRpWeLMtXFD+1wbtd82bBQtL/CCEjYUYwI8uFpPmoKJXdMYaaFbOJf9
J6gimwuz+SsSBW3Mb0MvYUN/7UVsP4JdZWdWalfL3rqLndLr76u4cEys6s2HuJD+
gCj6kurDy33gdo4i/4deVr/MTUvR3W2dpo1BJFkjiBxVvSxyPk6E2S2INUaF3I1Y
ScNc63fTlq6DYym9O1dbsl/W+EwvfLDocMIXGoERiDaQYYF6aLzYxv1UmzdpIl8y
nWEgz95Vle0zRy6x+Gy6lJKqPyDt4PYZGC8ZLaJhS5YsFPA+K9u6ZJSP9ATbNCSH
4lRRyTBjxRTn7fYMtLdu/78lXK96miaONkHJkFjQmjFUegIMueh+NVOqZ/rXkwkh
aD2P66OHqUgsiJyXGLux6mbeBm3kwdEjU3wN0mUvnyA5ZF/hQJSlJpWIobHTcU4K
jARyyoroE6wbaFm8OhRkPLE1E6dsMARzctDORwyeAFkHjS83RvZFwu92x4flAlBv
/7F8dVgwJfDO16ixYMWIOj6uc2JLTU62R5ku2XNnekSqOlpbgwRiJlq9mBj/Isfp
VnOyq2JuVsjAxW4SlrWNeNW4PwHsjAyOmzMwo+Gs21nEcqEWtbrrM83k3mUl7F7r
uqOaGQC4WeeKzemK5S/neoL4YQAcUm5F4WeSVVjN8HSShc4kUxO/OEGr6YRZyZtI
IWILlr1u+KNfcfGIGUzSWMpmHray6FZGwa+/KKKoVfcAAS1a2zQmQ2YfLgvC1zqj
daes+eTBetUzL07HhQ+EPkZHOA6lvLF5BG2StrCRz8+xblfT6jrPMsUbSt8BsRTh
WYxQC8PS7SZo9SNaIKue2lS/SptZXb3wh0005bKu2LOuta4w9Axm4TtlMUc8gQpN
CrmaLQcr77PgcAbmaAimRJNIcYazOhb/OACA+R9eLQ9Maexg1N4Po4pTEB0CbLsY
2h5yHwiTTAvGW2Nzyb5XB5Bp7/rNrUmRis71z/A2OwK9f53Hzyk8mRK9J4PaeQFz
eZgkkJAVh5av/UM7qkZat+H5YfFTEX3pFnKKUALmkjaTNU52GIYLMEkyYMoSv4gB
pwuxK/VUU9IObZ3pXcA6cdS6Vtr/wE0BROk5sy4bOB78M4i2sQyhXtqBOFWOBSEi
43Ag8S7jCz/v8/UPDBqdcE96+yf1oml8EUrrcwSyQvxR7Bs5UWNiaymkvKwbDHK+
PeFPvhx6b3CqC4PZxyO9f/UxPq9/yn/vUrwUWcgf23j4Kr3fnLjs0og+ybWbNGvJ
hfM63bB6hkcL0CPn/Z2Dl3i33OwQ5WpA2+I9xKZF+vz/72OaY6SPGPwPju1fI5HI
f6uVWetIwULKrWM7hNFjmhwZWXA9hwQwDUu05pAAOyWGBW2oGhzpaojA5iLSOARj
0jGW+iCMaQbt8hQqzsNj6XbYkU6RDHbrEi3+ff/lifqeITYbZO7Jf7IIjR+1IBGA
nPhjj9rIm9zfjdjAv6hkIJ1+fY71XMufgWqUKhR4hZfLEv9PGCKld8FNaO8Gh1Ah
CKOdc9hrUX+iSnfRmOiNSRpaR99EvrGLTgXICPDKKPXkHmMahlPL5fK4ZszFgq6f
XyymzXjnWM+kycUJXFkHYJkSbKolx/1ECVLEXfV+TVOuFb7CBsODXQVAg/6Z2Etg
H+/Kml3xEPMxeTUzdj0pgtBhQCh2IHbrKVp90lwX8VBPgksjLulIIfsdA0Roaxw8
8hq1lIpWgfIkCMxOurKafysq9SOG1vv1H3ZkN/Rgv5e0eQyzG7PTzSzdnKZKO06X
FoYXt52t9pv3jmYUTA7EFLM4GSOhN/LYeG2/uoLGUQca7NAt7I4u6GP8IxC5Qv18
Wi6ituLYXdaknNX60CYC5MmZnLWUuItIA28siPk7tQPM3Mux/DSOzzwWGWIp8L1g
2oilx/7m6tnjoupYzamKNU7q1aKBOUKirBLXdmNZa9zgClPwv2QCoWo+DvCtxoIW
fP8SMQepSuPodrvz+JKFowEEjPJx6TsMrXeSO2BlDP9wjoIMn11ESuLLwfvhX9v+
OgnGXZLsOzmiSNmvBSM6f2ha0dRaPMNEmNLCZCxbeQ4oQv0ZHGsz9od06a3IKxPi
W6ZbQmxWE8kzS1Su0I2nabkfnN+Hblxum1aN8C/h6lcemn3bWM4BPUprT5NYNC95
Sqb40oRVl6gW58/JegrvWAi+tgFOzPecAE0QYc2f603LJD1rB9vIHG0StHKs5HOh
W1yYRz1QZa7Q9g/5TkwsI11PNz6QIIGQIJgdtFKevDzwr8HkMIGE1/WecEaEuQU7
i3/XFVAkfq+v89eFgrL6PpyxhzCAtzfD00JWVGV8LuvG1mbr3hmLID+uwQjsZeOT
Bnfe4wHiyL+fCELPn2eZuXOZtj3cRWBkmpwsN3fdMIhlCIQ6hlkRPVLvft2CZDMP
JsN+nj4RN8V25xxV47p4cuE5huG8bwRAiTIjggPjtOyK3Qr+aQlGQ8ql1f3txo7x
dkt6iFs+ryh9RCDV8fdmN23H+kvL7yVGmkXmqtDqM3C/N2McRBxgRSIGlvbPfhDA
iwzrBa3tCK+KMr+p6nCGnC3gaeupkSvjq7BOzm1E04T+06ZeG5vn3qbSqB3frJ4H
BHcAzHz6wkKAzcoLWAfuwlfM4lYf60bhgMczXBnqrQ1XQ9zIwi6fkj1thiEXKYws
PYZ/1ERDb6PeFOZxUaIhcy/VUqYk3uaY7vHMGRii4dtipSsA32fsZ/S1pAyR1FgG
ANkVG+hZGB+eLMoOfFDkImNpL0xFkKkaWwd5ugPecokcCqeXxWh7OR8aZEhLpcFk
euOvUn5rKfwMZ91tIdZdAGuqQuNU+rldz42Zwg2XM/Ik/dA67DlMnzh8hPNzvwVf
ErJi+lf+RbKr3kF87d5yVriAFqYHjlSiA2IQLZmZSoQL53k1HrEjfjJlvmQSeUJ0
RSscPFTGzY6UO3J2E9GG3gbbTbG4nk2q6oyMLeeqwvd3oiNLLyao6dSkoo0DLgo8
StLgcWUPSzyO3goDVLsmk/a9oGjZk74AQTQeyv51etpxrXND6A8EQIX2+bUS8Pea
VypZBF+pqeXHBznq4rOiuBijt4/hThcG1Vi63SooqDf1mol6r/5KsD9TsyLbyUfl
/NdwMMMNPiR6cwUyh6IErkNvsGfIC+B+k2xLrMqJSgRStyVn5uoZIMa/WNAT8Jn/
h8MYAj0xdI05ojYuJiqq5qAq2NNhJe4UgzdzN2bbH7r9rkYVdDk4W09cerdItl6O
TYcsn55iRcAL44yaFHDmm3bcMcdzruj21qz679+flxXwGUHHphHMTMh28IEI0ZXU
6qSoBwpn9Oy22iWvSot5MHMJccn7AkTZGzH1ZLDJ79bcMB6NyETw064G8dXIKAAh
C9s4pcW6NROFzjy1jkxyNwVCGGTfBFEiEHVOBTxouDSXt3Hu3y6WY53KfXub+4LL
pC4kvEcTBVY4llOCJqeJfJ9LveLvXpADDuRot9oTP/uUDJ9+Myz0VyQqSdCA2eKK
D+f7zwenl825YZnl4wenSLnKqD0Cd6vxlkFmoub86tRrXefeXzNBQk3yG384gLma
0FNkFevkUnAIsKbC3pxp0QEdh0VjpCcAumDyIKWUmVA4WPaWPwedys+nHkf6ng8/
69CdI3GOc4HXvi4TC37HPwa6zjiZWqxde4iP2SOoOw6DcfVoOeiq7Sj1WDfK9fFE
hABqLaZPRXHBjx4e5/LgFWGBkS9nC1M8yHbiOywxWgE/Av3VyexcusFuZG99mLHU
OI3jylr+/z6KE8ZnVLQhgydkJDd4WZxymLaywF4hTzogbtPQjIMYPy32gXX+G00N
wxOmEVvDK2EKnHAqaHsmPetp8txYyn0+Tvz0wtikwrL2YDCdQ5dadvXWo1EhG456
HPgJRdrnDsM8dHSizSpnm1YjwtO7NJxoNM3xAV4OHPm3+mv+1H2FgijJ+2MrcEN1
vSggICz0frCJUFUNM9k34miAGJolrehtzC6KyqHZFFm8IQfCCDWmIHrxOjMpnpwS
2oagvu0SvH8GAkBwZei8gUZ/jxHYcY1j7Whysry1JfRtX/fYpILUrENiH/WPapM0
vfxmBiwv30UyIf3NoicaUTAcPBfCdeJ2TSPCOSwf36oInPc3snldSEwidTP9qv5r
h6fKSwp3B2vz8nRfHOnIL2KcX/2N1IC1fhU4usg5u6eruBqTYmCLw4hi8u/HdKxb
MsO/L2WbpGZSdM/jKufdc6sDdUdgcaCwKhbyDlSDdYJsf/y6l9Ii+I1QBU/nUjhz
tok3ZmSpgBDtE+h/C+c/gENvagxM/FmDE5CzOXiQGlwzwu2tFQ8tIEFTofMD0ZD6
1a6D4CB3hS9a/g7kOWNFwciJL2Rz15Si4IKWUKOU7qKgW2omwe5fpR9j72l/8tIS
kjlxEJ/Gu52VERQwa77wlipj3qGH8sesLhaqfnlzDzOQ3QU/rhxvyWRfJFicvDCy
PHGLV50IXM0mveteZNcf0XHM7W6ZqMXinzreJ/ocTtKcNDIuv5k+INSFLuUDhlwN
qb+z15l5zcV+qROxG57xP0oFsjO1rq4gr7bxvL5LT+55AH2WyZJzT+8iNNkhG0i5
OecVhE+lmYu2lp/yFuhcGGJldxUmQEmqUxQ6mcK6duOUitQQjaJJLt40Aq/0tl47
gGLvS9AUP0IYZJti/FKHc9McBw+qCuUTccxqODgjOpT+ggApNte2X+PxYF5OWmsh
o0Zvqyq+gEiCXBLF2FAQl/UmMBEGN1NlTvsVfxx14eJrGZuh25XS0rNZRV/VpeFp
e8IeYswe5G6hmpoXb7N/m5+67Xi/GURy1zbejM1pjNRHSkfhgiFpEZBWthhEGfkd
rcQbmFTxEaEZ1NPPAkWQktvu3kYRDcrn/NjuAl9V6ME+QAHj4o1xNAX9ZE9q9IRc
TwbO2cX9bRFxQGBMFDB7MtgmK7/sr+gl4lK/SRLN4qZg+53Ti/DB4+8gtwe/C1Ic
9Nt54n3ipx+2jEE6iRdc8fgAjTWUTBf6tldhYr1LWWb7uczr1oW73igmjsd/GnkK
4IevyrMk91VFXARoWCJXp00L2d51oxPiUw8pNcJxBwGQKSylvvyBtq6tbC983pad
zpta+BXkjS4loTtN3LCXiY1DGjQy98COZqmkAn1H8bFLtspHaAna/mDASvQ2qWYE
O0aoe3EFktADMa+N7U7e659M6Mn+DLvfCsjlvcg2/u2PZ5c67o16wAv1uI5pOf3N
lGoHfqBFkLmOrGlx+LaHL8Q54sGtQ3nJZAwPqeU+6Z8hc11vvNcbj6Dj0IYrg2Vo
Vub3VrF43k8tw/MUsRwakpBHU32evZ1CaIahQm1ZWyPBxXhzeVLaSM2aUNlga5Nh
lp8xZAOPnStJLYTz3wmiPOiiZl1BND/sPsqIpr45YYX0vIrlPVg6tjssxbvamIFN
5fdnQSl1Y6yCRbh1ecQ4YsivNEb0Gbn4zrtsA7L0nrtqgz2aRSydPCbssoX/XlA3
hfaiSGyTQQ1fiPsPRit1S9W9CjWtM4VZK9q+i08c3uKQ+QBkCN1C07cEmzTls029
u2iHNT2pgL2dV6bvJclfSuTOBY/adPgyKUrpwf0j7RTwUxsDTV71uDXU6ClbI7xU
IvuJ72tSyR+Gg9y2p2KuZWxq8loijTtMbUdTsbkAimrG5IjHDqHRbWWimkuVMZMs
Pz04IFrAIgCuL998sXR8k017aSrsbK1lmvT4gRtsTpOtdRkqLjEM3HUzAKQ/aGB0
9eGDZWV5zv/TVLlV0qt20DVzKIrzmWvf/Mo+6YJI79lWUbxnoVfmtcTadV3UrYFJ
YLJ1dMBKonFeys9MNxlEKd9kcnzErxH0KYOJQFBzmSTKXUZcukLuuP2+s1Z3wJC+
g9X6vfGXF09yN8GF7TUBBxa0tnf0LnmT8LF3GLk3oNCXME6yZSX23Cos8B01cGTu
9lluMjy0y0eLYKjrXCBkqDM7tHtWuKBUAWI1K2HFdc+2gqHmu3miTWwUAmhLszsT
CCPoH+vFzqzA+OkXtrn77uqC0kklahzyoVy0nbHLVhPb1r76SJXOVw/ioZ6L4+/E
Cmmo4eLTDsTdcO4gYMeSwVsQa5rIDMAb9tzVnA3BctwCMUCFfx9yvvis3MR3VRvh
fF7LIT41268j/fzmnFF/M6sdxAjmQ7FBRcPuAYHkB0XRsFAUvgHvzUnLKYm+LniE
jnx099zzwq7z/Uilu6uCgFanbz2XKHn+OvWeBssMiwcnkHSsbW5+A2jjM16nOfMl
yJiA/TCz8nHMBU853UMPazN2BeqwFrWdC4Z5Gw0dP+9XH14ADNxow5t5Cujq91Ba
Wt4ONqKAloTtR6j4bFWO8QJQ+NQHsRZC7cd2Qe/SCsgs2B02ZQwEfuKmXSwl21Z0
kc3MdK/fFMQrW5vYQWUfDS8boxRtCxminqvhbQkI1mswd8avDK9gg2gltIwVM6XV
dRKmiJM6L3INb4IgSBipnD1gbkgH1+4bpy7Ld+uOTmm0L0Cv/QWcv0DfMjm+ZDXv
tZtAHasFVdv8gqJMlYDH8FsV0kf3TgNktvllQfBOFiP8uSUr0F1TGJrMrxvrZrjD
pUXoBpAeB/MPUfM36cSZ3r4SDYLVTSv5dgeSXQU61wJ5q2zthbyd2LSvwIi4kTKz
otMHp3fcTvmtRPxfs9DleQPpQwSSgJkgdaBKTqYup3+W4UoOiMELQ+P2GY00dJ9+
XAxAsIej5dkdNyMqtPrWdFH5G+mFqMDa685XytXw5h5bYYHGTxB+G6bcPBAwYd86
1Dtirmduc/Q4da15Uf0WJtZCrGeA1eCWaY/XOz7ltfO3XmDt0Do5g34PBTUTYuEZ
ztsNrRsNPC4ZBd9eRw7sbny2KFDK0evF+UWimGuUZcb9lNNGeP895K2VOJZzflI+
yp8G+PUOH1TvVdNatwQ9NeubBIiywh/DbsvYd7y0IZsN/QDYTvYsNUb/zYHPGeUQ
bLREAZRWFXlMYzTe+P2dnsI/r7hJ+/CXbzV+FeYazJKUrU3iy/bmzkpMj9EXkmHB
kblp57SZ4BS4DLE6NvHmgyua+Pt9P1M8o62j+tI3ypf9gZf5g0vtBTxTeTC5nbJd
YpSdVowButngWCw3H44pwxYQz2TuR+endSg44Rhv4UlJh+KCdBfTIpRE3i/bkNMS
oYWANGWDeu/WQGcl/Ykn5y+VBPgIQIOtV88Ky8Udssih32lma7GbLjoZ47pJcZX8
ClTNBfwcmw3avjHwiegbxvHNTEyC6fQJBLnu8xssHA8rF+C28lbpSOugBlZAAVpN
rvU4nD4lGcY9j278s5RwQeE7aI1CN7sEt+q6l2JkNHuJFZM+GH6pjHwEF0oxIdPm
dtpKVLJKg3c4shAQP2o4ar+K7/ROm16jJUTMzPhJYds7xbyb43Z8RbSBAMsofu74
tCTvrT54R8EXgeNWaBd4QDREoVyo4Nsx4mBGe+tvUpa806zVN0NJ3sC1UmHK00Br
Fe7+SqN+Y9NOOykfrBJs82g+6aZnKxiLZ6FTJqK0Cy+MZN96HxMo9rjGR6xaiRK+
Lz4LpAyoZywpBDFSIMgwT9TGraj9yt0WAgOxCHv97tLC4M4bY1EMlvINfb5Vq3cP
3869WqU9zm11BqfJBOa0MZYP2/s4EADgV/oJN2UtJr7dn+PP4zwAvdJknEtWYblQ
FKxt2Ffwn4B8x3v7Oct6N1kyc9+JTMe5Ouv50XBajBMR6or9Wmom/LS5e9lAKKrP
D0jxilzRBf9V/wY9e+4iB135UlVzUBe4epgFAsygIjMgQJB4IwCqX7XKh53iWZee
BIeCk7im+oHzPfXS/Rfx5ijtA41jhYAtqz2l2FM3Q+vBWUy7RzGjwEXjgsxUcJ8l
rIDh5kGLONp/Hs8r5AWP7Clm0BU0pgG+awvUs7vYWPMAvHDdQkGtdv93OxsrMX8U
9wCKlzqcRfRp5sv+/icMTcZziquG456IAvRBXN56l5hLargGiv1cfjv60pswNfDB
vcg1NIHwfMbXI3qTihQpV/EZ+Q6idgltY4+PBkUcNhJyuqjPYUF6f8p7+9+vc2uq
CHFhJvDZbdkMX07J/s9oRMjJw95Cyg9pP+AG8lBxw9ARCyTWd97tMygXdISSpVyv
DYrteEEnHeQ6QX3qcw1SyYb3suWiYTuee/j2UUtU54AEoWkRLSlo435zH/R7e+Ks
0+GOPfTb2tWzF/XmaWOK9S24jL6OQf65wiZqheBYVQ/yWMhp4EBpsQvV8iR6ahVm
n3XcRmFBq526++QJF7alEfaTTiJkhrRPqu4dc31/zAs/Kbj7+icIBRdMVol+/x98
BJwhoyDqu6Osu0onFHrMuSTi7ca09yTQxRad6ObhL+TPmZCAaG0nrmleYPEP93tD
gBglQ8vIwJkY2bCP5aKxBiCd4zUz/23SZNvtwOgm+8cMeRZ7y5DdM2ASwPDA013P
yXIjJq6BlOyXn/j0px3+EMFgc4FYyoALBc1PgRUrmr7nbNCAFj0wPykih0RTBIDA
lG4hLtVGkCumDw+/R1nwPF5gJcLTPLFuc9ggkO7P0cXTEHco7vd3Kw54UjYeBut5
Ho3T+fjIyZn0NuKpp2gfm1jBzlNme8mLxl2kBMARXrUEQSF7tSOGLe1jm5IbwRTj
ut/TAH3nD1IysyDyseUpdkrDVCCOW4Ryd1+WoVBE25URVRCqtiN5c8IkQdT/tP1U
VfbJaz4zdFaFnXgjhCJvmz42oahc1/o7k6uf3PffYfG6vU5cKUmueHNsEMV+54O2
piIGr+C0nGF07u436HCne1NSTSsTopCsduQH46/gWdBGPu7I2F1UXk6CpdsrNXHt
30pBLBGqJ9hjn0JhH2MHCnx9E0EEEGLjoExbZ+7vWNinDyc48Z/CBHYYx3pX3aOe
8h3ASOoZXeyBKgl+T4MxjbrsuBR4R8PsGnfKhKbUCKyAC9N3rUFoh540cpFojtIi
lHfe3yL1qnG8zqQlsCONLMzoXFY2tZxQfL09O+HFhHVLIdIWDKr5ybEwLbbPzw4r
pnYElqgwH/v89hyEhtx/Mp0t8qLZkMaLkYioIYmofCZ1lrXDikoutbhT67PUIp+r
1CcN9Z0e1UfVyHkB+hxgr6+a0Rl9KqUl2uRzVez5vjzrwIhFoZ36NJ6VOAkC1JPy
/WUVu4xb2qDDHOXFJCrvFxtCSJ+AaDHUrw7vGDXIO9OVYlVMVvpRk2hZUcUR/b8R
Tx9sLnKjMgAjS2Mzusoj1ZFPPG+8QX8vxsu6IXSaO/GG6ZaeiMWjwVyH1uWe/DQn
jR57j28Z12+Nw5GHdlmW9fGKY8dMrSzm5CTPSX40o+q6yRXmMFXwh/4LDFA/dkEo
wtW5eOHKupwWZ8ysj9cH3BaB7mXMjvSUvoDQa8oA01Lihq1vnzlHbYpjLZLont4S
NJAATaZ8/EII58zWT37pgY2+6unlix/kuO44DPcpfY0stuj3CEOlmQ0EGeA9Uqnc
wh30hOYh13bS+Vnm/UzIs6vqqr2yHAJxV49UNyNon7oVbsoNnwn4GmgqDsSESPm4
ZNxVpmGby0yD8N78kIzNw5SwLoB0RMm/1ONJG8SFGtI88AwbiKR0WulUCqE35h7R
jIzPPYjUrgDM6FTznSWc3QSNEzpQ1wAmprX8SEKf496njX4wT9fAVteXfuZ3Prri
bUXWN8gikj/mnwJ3gPyqbfnRIHh3un6O/t65nZS+dKgbr5RAfwrmN6Iua99du4R/
U3iAFOY18fQnnzDDeR+8jOEp7h3pz1nPdWB45GJ1WsOTDAyIeOATSD1/QxcRe0rL
DTyr9IwmY6Fokzt81odMX3ug4Jj2ZtucBqrLmSl/rImzN3WpnKpj8LmDAbocWYGo
wsZ4qJbLxMzE/6vcCFbtj+zld0Orf732BxMccI4uUzyA0U9XPQqu/pEIkRSNZLV7
+pWPzENqDAUQvPZIPobYlHreVEeoAqfpyvtNVhcEPzVNdO/hZpvbd3c84QSRIi80
UfAIG4WJIE7ZwD1N5U/P6CRQ/BQBZ/NKCOK0HkSeQ9KIM6jJOmPayO64dLUlsuEh
fqRnfz5paRc0EUWojk5A3MbaIwq1aONgN+jiuuQ7CqkcQnznTu9dk7/siCdCbCas
kOT8od/VuFKncjBK+ngoLKVFArlk7/oN2lbieS6j39LTUNAKhGYmrCw7tTwj2JDx
49RCtjyT/QV5FNQtsW4/uTHozLoq/yU7WReS6KEMIUnDAArBqYfDTneJV/gZdWOX
bswBCfm3zkhrr0ZY2b0jNZZt+wiuhu1G3IAr084+F18QpCOkxRJ3nScg8fpRpYjv
wwf6QTCkNAX11bIM3oyqjgpBd0IRIKBWnzeW3k1JZEinA6bdt/HP7Y4AQe92vOeJ
5Mx/gKdUR97K8z37Bz52LJk7x/RIoIBa+N8YTYP+3ZHZcPgn+KIjdINPVVBfpkSQ
LZFrBG5GSsJ6fuHjEoDQWwnlc278NyDKUj4wv7iS+guJJ3zHYAl7jn3CpPNZuROC
4Oo38mOtX+snMoS0BNSvEv4iBxl6mJkKf95J8pnqYb/kHZJnATftHplG8OWY3y85
HK0RXD8gKVe2ngs3FIDHp8nvJ9NB9OaQ24uxzxSdFY/mxmhq7/meARYP59/yCp71
ONmNhbcMiNyFAMFovghWG56tlqqm/tkd6HXCmE7FMApwinNNe5/JIpHnrpi3xrYO
F0Ao48KeZHMKeeIkhkq4NqNhQXWD6xbEui1ljQGJNWP1NpsbGnpq4xLNF/CJePxt
OAeO7YHBdH/j5CnNszkK2Fo2zXuQlWwmB2rw/nT/grjvju5xSNWAytAHlWOUL9MX
hVKL0s0QS2Ro2Q8Fzh8JOLdNRcoufD0OSKABXK7f5A7Kjm/ldkrbXDgrnyyyJKkj
OX+7rtBpPjBncXVDxoZGvxmX5q/Bj0vdBbYFrbs1UVfwIMTgIQ/kO1uTEZ4AKnBV
6lQcjS23eMGQ4nOlyi6rKNmGgkqyPu4rGuBNA8crmttBDQt1q5deO1oF8UeqkGym
MQfkkkh9M/Vv0ywLAS0Fl5aS8N+JYizA9HB7hn44c2gTTxzy35EEHsoBRsPNkk/G
dmmWMadvYhcOGW+GT3fS8Cn6ugAMt5DIrD2GlCWeUc0BMzqXc7/Hwr9o3N2uO137
AFKPPzK8vpLDPVrPYLqQLw0wGNZC5bnd53Pl3ND3f08Gt8tHKrxoqD+u2baNywZE
+Vz6g6wd6VLgKptz9odU+bIz6U+baVmoFRvOdmiUkjE+jJFRN9vbbN94x9T4HTjW
ax9pSWk8OxrtS4TaEui6UUGv8IOCfXvvG1kUZZ1qINofaZ3LLVjQcUuv8MTuO3uN
K/Rw5vANax8WW0zQZLEY/XTAsXFB7oviPpViEX3yGeTwXN8vzmZsjgDAwmSbjULo
hVgtLfJE2x5z1piL1oZg7K2cJqQFHQDcr2hBk4+Mj9dVJf8EJ1USilhRcUk2Z8Oy
xdya8wHtj4Y082ySGsao/dWRsa+hiUiLrF5QB0T1plQR2KW/COMH0ZmUYryAqJ1+
Ce28uO52Kvhwseozt1/wJbs2h6pxWPGukIIqmeXOPxU1iMMah6wdok2TrDvZc0eu
fYplE9GMjpml21JH7Y+pVh7zKKrZQ8YG313WSLFw433eynVLcuEgJI0P7+pVd2rL
8tHKoZzW2jj6oSbVD0pJP897erNsJelZMe6hComNGmfyUDECmpgADljWokJ9wN/t
DDmbf1mCfzk8rIermrskr1X7YRAndVguCQ9+WW4LJKCpZM2JDGm7BYKZJJROYaAT
BBw1MeAc08+aRDEGVY9WPgv0vskgYbUIqkbGO0av4A3ZCFZqYBW7dqwMI16ioixB
B2l4ygWVemYGEWDK1fVBjGVW96WnU2HhCy/hRAVthle+/TnPQ5CY7XN9vdCdrwFf
uojtvylknZBTqP41hUnpM1I8fdlKK+FOszKU3xKCj2uHs02oY32VgS4+ocnnZOgh
QEnqCHGJ1Wt45GhWhFA5tfa7b3jbn2HyAPDb136EN80IsmWsCsO2d2cbcr4SCMYI
Q93zVrP+QRLL/2udfulydtpkzXAhbvNUAMZHFRI6vptC+vxdT3yhmwcSp3uGNH8D
w1HeqW1iuDbAa5VDK/Xe7cUIOuOrnGW1Jkh1UPkqUhO1qWhO6FfJJMMDEcTGgJdc
I81uCAlDUl+RsEOUv6JxUzt7LJsE5cV8S2I+ZLCKQW8DOZEsuUyvbCNEViyAsmOm
FYVuiXe9+JN9nQCpXyRdRwuK5xwbbpYKe5X0z4jkDZtyDQUdPlXWTGBwtTusxFP1
jItXG2GDD00J8zPTChpw011tDQsbYj4NI+a4KYsz9Q49bKapWXHFtcaKu8HYJ9JD
9HUU98JAzusBt0Kgk6p1hC87Plpkc4DlHSv/pekfSiXnf2cD9ncKVdMbKcYsNMBf
7vQb9VXWIT0dSCfDIoOVELjuFCWQlFzJ5G9dzQv+NnwPG1ILdBy9Qi3JAlJjVaxD
TT9ComJitzK8qkYMvNuzvXLBY5Qcfqd3sSVWgjPDcw9vcDRGs3nvTzv0TbeHA2dW
RsKMhD3zfRA2bL5lO0qkepRp9UN0/UaFd8rFm0RR7BYOiklzxCNKO9DvpDaB8bhI
d/cXVEWQiawkZtBhwCgTazqe5TLGbKiUg+IyHN6UiCjw01oJKF2WbpaB+8UpvBH3
+S9jQItqgwBvM22uPumTZoyOV5eLGJ+jym4RC+Duem8CGMXz1N3laioaMshXrKE/
KmNnxsFWPeQ97kFSePj3TJ1DW0ygdbXOdG/LbgWXGbet+Mx6Q91R18jKYkgJnaSt
rL8E16Xx0vu2txniqI0/AvBUAC2snoMyeNTe9nMIlnPuUiOJdEQMglq6Tp4R7TZb
s+tm3Z5DK3jpTx8LVGmlOW8eLLmMfOIxL1HSvNMD0hMN8rdyZfnaWRrhghuwrW6J
lCUB47DwOrkZmGnOBMMR9CBqqLz1S1egbmL2NxVu7PdNzV9TJB6CX+K2NHCMxKV7
rP0cOO19a3i5Vz8fF9xDdecsRJwAPfUatfP8VnlQg+ViZf9dSRpjha0pxe5pL+7C
wkA1jhi2VwwtQ+QoxCJ6soRsPjk7TZqiP4z8VhokCmExm3c8YKsHAaEN8O96VFnQ
jJz+m/edG6V6xP8quDEcnBhMIPqGkKyMQasGupQOZUZp/u5bLtx1iA4OspjxEVVm
2j89NirBGMCl4zRGIL1qT8+XH5M1EueM4CoxXsbfACyZQSdOYDaSQnj1j//qDnu0
VAHqANGjt/pE64P2e4iBsCOUsjPzEWPhVfF5kOxXx2L4cyd+cNKcNgjGUXGKOMCZ
uq03+tPgcc6I/QkvtzoqsNUv2muuY7Nc8d5hjta5yY/w8a9bYz292TBEKtgZJzQO
QaYnnsJVEDTQTICNPv9lshsLxVJhqSxJquntvwsi/eHDTO9HWk2/meekbg1n3G7t
v7UqUZyDK46F72QATgy/r9MnrFc8KLInLfKcqPXeNzsIjmcpbhefUFLxEKnEsKhu
x4+oDuhLCiX/eJyY3DfdaR3/EMb3hrYAuXTU+8q1Kd89Oa2ub2ag5af7IyYQ6z4+
FajurKBeJ4pO6Jy/ic0lpQL8JviFySAU5MyNgGjBcNlmfMIkWiyhmfGY9rhuMvvC
QDr3J04r91ZweS1GqpTCkRHSkrrU1doUOF3GJ2LqeUKwU5WgcDtepJB5gwbjVKfV
U/dXtkq4iD6+TLgSzgfozmEqv7zxGTSqDjtWepZ0U3ja6s9h1/wJqNz2EM6RNQ9A
50ATiDJRXOBo9/0C/vQ+Od1XpB/z3kPW7/OyVHxPotCF6IFOYUB9Nt8m5n6j3BCO
7HbDbf9OJbIwlR3JdFJ5e1vuAtbzgJoXnuSFNN+uUpMRt5obb9Pu/bNHjQWt0hhi
TGf3pjx3thS6vIFx8BkCEw8qs8pgGXetAwVGm9deqL9KXdJc+aOX4+j6xtwYzGao
C0iwxrWVfjf7uydg9W4pj+BemO2aAE38SGpjpqwWbozvzVew5YpAdaG6edmLx+0P
qvd/FkT38xbTjutr+BwmJA7yHV9CYeqZmeCJbyHFMYoi78EL4Jy+/NuTYUUTMvbD
JfMe2btqBOUFJoMx8QyzKVV2kQAvIvY5g2vpvWqAK5nwvX7flCCn0WTSne6P86lL
VH7Zn8iQVsGxJMjwdxgKxIj3ZjE372chiXz41g6vuKfzC5wOVe9BjS+DlHtR9Kg/
ZJrlqJyhk3DPP+5uNFgmDHPmJ/qw2ZaYkWGI/hI+a+e5zRdi2Rv2WY3HHfi3Ky1F
cmFpjpDz03Qdo7GWja1lBqM8U0feYcQxv4lBu1KfkrUijIGI/wbFBrTLg0gRi2cH
Uzut0Ohw/4baobcS/eq8lC7TjoRZFkU6VbgtKtcksVQcj5MUnIIaMyqj58H20tvm
0fRyFP3TO/rVAIzwafH68GrCC03+aJBQjnYSwDAgj877LQxp5sOfybPM+IAh7wmx
DtHlgxAS7fEIzk3ESrjBpNLcUFgwuopgBrYLV1zy0/qJ8+fY3DG828NB/SzvuRFU
hsTYyO+x/XSc2xONuQU+6FUG9eq/R0yqu38AfhtC952zH3wtwejBJSbYNjz0le1z
nWgIeol99nnBZcXniLmtUoHwLI4i8ILPAmDuVGDAGWWLe0yK2drNEVRkxTGiVx8O
yWSaFkySs9pCVCUXyNcUA/MAq2wk+YpGHz9J5S6xGFvMfP9tsfAQp+ONef7c4g1d
SlJWleaPeX9HXtMAT1opAXQ8r2x67/kjhus+n/A8XJ+UnV1fu/+5CGinAEUpwhA0
N24WBK508uwFgRMAxFIb87y0pCM8WoToh0WPoR5Vs7fnE0ogyH5PNxki+wYpeLRL
9kt58Js6HPtwnYFDEt4ggl6rmhceZoLKJ1yZUee5rrad3VjfTW6YfnxgHvdkUvbB
O0dSaU5Sm8TZI88L0mFg21nLnik7cMb2dBb3pGH4TAhas5souIc95dClUoLUygPX
YrEjuJFCgOcO3r3IPd6coOngQwyi8JJs9DpTdjijq5oLtLRfiVRIGSck2U/ifwm8
fJgepfKflz1gxdoh9UE+kouN3MI3OwkIZ8uDd9FpA0e2Ij56R4C+vGBVKwkUUEZN
hL7IHZHs0jeAB+1OrlniO7oe9dw3w5dC9inDY7u6/beSvOuG8tDfUWLt9o+NBPXx
uEQDPAswtycWN9h7ONvBnEDFemK7ZesNtWS4acR52XCntO3n23v4vrK7e3J0Gc6n
bAmzETeBv764g8BM4DA4ZDik5SReBfvUZVMrMvu2n2e7+8o+zHwJQJhXujcIfgie
yS+2cbR3ElIOm57ARP2c8nO5113amX4iEG37p34U4ydBmJYIv3yIOKAGtSkKQb7M
rG3HQtchpKwiZXk3QoW6iOWDSVffG1rcbGzYnBgJglq1QPT5/Y/MOwCPO04NrItF
WjmUysltjuMHqmqOjVB+mimmPmKhJkxvRxyxfhKeOu/+OY7B9NkKTy6P/6sAoly0
4NjYWK5FYtoq8oLQsG9Lme9pboXpBWZLHkswLum4Fsl5VtLc3IZnqNyA1cWrpqbN
0N/re5LECxN9ccBPotfNRK5gjhn6vV7uBanQk6Qo6/TcatXXIV1lDvk51ZqQPPMt
HHg5MMgp8HGtw6gmi6X/HuS7V/vReOZQTPvZ/5AZZWsRJwQIVKTZU9RnqA7K9HA7
TrCPMNBsDlWH+HnATqWFO//eTbSlxg4pyr1F7u2iRaLTPsMffXOr8vVi6qNXUSGU
PoDqClTd7zwg9Z8Rp/T9ji2Ins5tL/pnePnzhC5fjPOsRz+PZk86/kCoI6OYnAjt
qVMB44BjEP/FleG4hlioAsPRLris8QYLXq3AaAX4gAwUH/5/YBZ9JmJ2f2Q0ysnw
RjWqbB5lpAitYGPJX0cVaVq9XY2gXsLyb/CLoB4a7QYwvVIrlQshwN0bIqXQNfmn
YF93hWEI7G8HJRtLU5dRpVX1pXZPUeCEbtFsFAY15XfqqsG4W8oKEL8CQICjRVkd
EwtntIdB3fL11NOYmAMRkFTEevJ3QLPMfbZeKvoJLMMhJM0BD+cZZXie+wgFqg3t
0UZDvm03sCE+mKDI9pU3dLXxN9uFn4N+v5LIyblstQM1G2zGFX5jsxarwupsCnT1
vj3qp4KG+goYoNHM7MZ+SeNJsrmtxqlNZ89IqY0lwv6vYaUX94WrYCfc2fPu9dZ6
Xzi95Hm0qWZz1X98WRq1VQnVK8VfzPiEQdTAHHl796975A4Td22+IcSu58vWs8db
15DcoppDeVFX2mEvG0AI0c8K752lxFVaYE9Ee9AVcSWczSgLtCj3eqAzTJcY9H+7
TA0xKSuZ/2T3d4cc8/GU6VnpFcltKovNKWN8I4QrIFSkduI4+mQVVho6bS/OGdrm
1KBFm7ltVwZBHQNFqI/mKN5qKw6ekVxUpTA7IVOlrVz1wvcKjo4aLubdAuOymGcC
xhl2KqvuPxNv+FB9/May8Vpzp5ArXgyjvsqqF9RkRVQ1mPlgB7POo5Z7M101I5Fj
m6gpgQCm97IEGi6uOHyXtb7L7omMNGf1tGruSur6PkEc78eJfFLxSJa1bpwHtOL4
Hayt5cvvRSwMzFuTsWEPK9SycZlNehtUmn6mo4hApzxYuNkBL3+ZzyzIH93IkhNN
ucbciuvLvxrtuKBztNpIrg2Uq2GaTu8mIPouwwmtNvDQYIT/bXgrR5F2xHkZotwW
2RANW7fBy6BE5QEmhKUx+NDwJvYHGeVDRurIsm2Q9+GBExafLOwtf7vV/QOic3tf
dla24vCAt+UdZiYnpyKp7cIXB4drsGCxhy9Or1tHGwDMKIBQWsYReTgLoifqgW8u
PfqE67isdshahvbMcMSy2XX86OJ9B5zXswN403UVo1cx6/A76gLLzOkHBQpuUHZ7
menovDJd+64gLTaesU6Llv/6PRqhQJA8i4iYvyLS2CgZB6JOKpfjSgh9N/OvIj0P
Fhd6hb7//8d92sWeps542/qqWYka6VEwYPoktq8PcsV5re3mYABWYRyYrt/w0Z10
v/miCidpOkYZqdUrE/IaSXdri35qD2bFU2c7B5yQOwEJ/dBVKGdIhAnLO2pKZkTA
048kvNfk0xiT/p0LqwBDWEV3yQbFC20PeJOpItYqXdfvl0nIeMGgAUhi15nTfpzA
VSOcw/mvcAJszumT3zsBCMIaqaBAcMN0PDpCii9h1w2tR2ilcGMjVWIV6QQXA6yS
ndedGmfL7upiFDlZt234fiIn3zQC9V+VXP18yI4pGA11fXsBBvij+nV4UFRosd2G
QcPR9TZ05ihxCWjnUz9Ej4p27CWNlF/Sji4/8a8ZeXrwMZhkHgdfVHa6tklTl1ld
FWIOK7SGgeSpQLxCyX9Pn8Ep/9EZfZ1wS41AgT1Z/D3xknH6JTVocQMmlXZ3a8Xk
eqrawSSo+4S8YAOyydxZheVREK7XFZJzjs/IY99vUBMWCDtbkwa8+ftYvQkqeKBh
afA4WerMn6oOl0oETwk0jkpouqKSmFvA4KDKPK377lhRIwdnNwHVUvejBKpRYZpw
Vfoe3flaHDVEv76w0ue0DEWVI6chxvBhtdH8spONDru0y8HlJ27YBcCkOJThVSvV
0PZd4hlbyxPrvW54hMyz4vUEByoFCMPJ1d1hQkGqKRXXX/Zu68/1LOwHoH1259GL
sEJjGNz51H2IbEZISOKuf3jX5AiMk7tvL8UX47K+0c6A0kuyyrwAmupGZsPXltRn
5T2xQq0KK0m2C9Jarhp6Sc6LK8Dpu+sHWQSWpFbJ9JL3gQ5tph0at6BMNg+FQFOg
RB92W1QY8w/kxkWhXc1v+rXeQRHZSrg+BoWuDZOkSXs1wr7dnCoNt9QWtcpuf5RE
197eKUxAOUTc6stwyblUsqdUsmVz2IwT57tuv9Vq4T0XwzASGpwsJUdvnn4I1WAz
mO5w6nN2KaCz/ssqRs3SIaOMebwbObqWurqrpAfD73Nl6RB9dmg3zDo8/0x0jLX0
mBDEuGt/5vArmULAEkEq3qMpqo7NpLB3vHv6oMkQOy31cEQ1ilnzIl464FmSW8/n
AWwgkEsUFYlIBTlePQssz9imStEpSwnrguaLHerl1gUC6dmVZaho1vfTjJrV13qi
nB7wZ1xxkkCDxoygCl4cv9z6YPwbBYuDzzASWIHWP75FRFeQ45UiCnWMc2XjHFuw
7yqBxS2IBl4t9M6oFGMqV7beKK/YbCNZONc6xwhmq0xJXb5G0l53UN+70ib9t7c7
eM5E7V9+wwyfsvIE/kD24WmM1A8ZEQYfZCeagQDot8LyW8XmFFSZJysOQratfAkV
CaVzUzkEi1CE8HsaZNDwJQY911PFOPVX1ltM5scR6sq+YL0piOJYTdslG1REj+FG
VGF1lncz2RnlK9xTDbNz07zzqbv8P82GumHGgTh1j0FQRl7H1GLaLOJ7AO9OdmW+
HaTg1JjV5inBTaNVFncGEwpYLiAk127zxsh+uam/tbJ0UaHsXr1YJkqM0dLInjxM
B1KvrQjXeM+j2hr5pwG1W6UPS8agrngueVbY2HPPZ691JXrSp/qxqV4LlO9R2hKB
Qk79gBb6UrfFEOZeoXZZu2ZmILTDSr/SJEDkfu6UFgi+uwIPHmybTZvpTk7DXMlZ
m0CZr9D1OEnTXI+OuC8rDs7RhkK3Ene3IrHBA3qzX4NOs2tbsCHDEYNVXr8g6Hsw
LqFnkCkix9IQRV35ePKxsZqAZ3HFQif7JoBK4BEUySaEVLbD/IASR4lAmcMGmEeO
RjJTQbrjf/u2Oj/G6zMcfSqiWvtqwd452O+8xHlavH3GDcZP4LOyWJhux9bXSj5x
WfRQDH5uP6LFFbuqzMODCOPyAr08OagnFlSTKY5DLJ9alxDN6L4THZMSQoTfrsLQ
Rdt3Yvyaz6dW+B1ks+Xf5ufWWRI16TAYkicESNGKdhuONeqIYv+RWZCD4nkKKIsY
05Hxp+ffa/t7uTJyNpcEgx+pIOtJ4wZ+y3lP/LEHyHVUsFz64hzt3oxJb7NSpcem
KBUO1bj9kjf+wT/CWv4mDy/P3exX1FJOz1z/5onRv+WcAAC/EAzv8kF67wr1I6fM
u6b0XMSXefbkrTnCOD3/cWE5EOnXMLf1na7Tqp9Japkm/pfuZwdGlHCwrlrkejQP
zrCGcPff3Oy/nTVa+6jAdRqXBM2ljd+hmxNJK43hUtge+q94VAkAcvRzwjdkkNHA
1IjKLNM3fDGhdAIpKspJ6bg8OOeh8CLkjH7rCgP+gQGV1wJkfs57zVELRmME//wy
N5nnr7Nr7nQ56pUCD3fSwqvC7IA5gBjpOR0yVlj1JPOJe5ej7XeUW2sTfa6RT6dB
K1P6/qoxaA3bkt7J8hsyQX6uXKRVvNI7VLoHmI++Wtm8a80UXCc6Oe9tLfRnZ5Pt
FJdjfHB5X1lRCIBp3Vv1ne1YU0/FfF+wFb4txG3W3gRmnAM55xubhvNqZq8AjrZx
JPRsESAuPGSkhGmg27NjWLiaX+WRYOZ4sBc8UKCL/F9ibce+F+/5G6nM1xBzytfy
sisAO7hSDRJZYOSzy4o+/6QW/cjBOwsSrq08oFxGuDAxdINEugVcSpOFf/nZhJFP
UWcRO5PMlYVtujbaTGHzpLh0j0n2jR3OcNQTOyDeG8axy0weYv311ie58ufjayrw
ZSlzo76OuApJrBWpKijfc6aOh48+BElX+ENcker9vxWorDsg3sZouejB2rsrZYhw
f7OrgJdBzQb/eJ+Lgd8aNQzug4NRWfmuuTi+DXoxtJCZ85+kOyuC2IK4RNPEGsLC
smKHGKN7CRv+ugbToS4QtZbHUv7nxC++Kkt6+eb4wEqa1C6Ku1PHEZlMA6SvwFQk
tE0RHrJHqbRX0NHawHv8QDlv13s+35y4Ko3UMFT1JNMoGsZVlxdVRuwZ/g+/u7R/
3IHuxQ8PfE7V9Z2GApFh9EjWW1b9oG95PkEeVZ2AZSTL/58LERWRWuIqj4mAviFM
5nOBWrA297Rlk7RxSqcsB2eTUtwwTxIKeig1JMC9YtB0ygzYGLfCIleJWzcBCL3e
wApu92gYEZg0CH0aegRP+dAaD64yfH4NdeTvMPfRAoZsQGf8jD0Oz6A6y2AePjGb
2dtNxniFdfYrEupYrjxNKt6MDR3+w0ElC5He4L1yM/gss5FeQDC5529onJEsiDY2
cV7PmzT9FI/FgDsCEuo4DeBGvxeUpkjWanaLRb8tEaxxJBOXlWi1RuPxdJAohLjl
4ujMr5zef0TfWUKwTnb/6kVWaoaHYVLnvWoeE5y6TQbVcu4PNa9mIKxPaCu9RQXe
KJ4WBS3lIT/EqWCqDHXKsNpgMcl+Svw12K8Hk8Atlv6SpSeo+eSAfP7kLeRPJWCS
BQ0b3tKjcEWYMpb/OyQROYgqEQAVuH3JZ4m8v8Ez5429ol3opFs9uTd5c7POG6hF
zUgd82xASur84cMXtf1C6Wi/451qGQcy4kbery1VLeWVDJe6Eu9X2O+NH00ajPIy
N7mVnbdmYSoqYMen3SclYckQ3DJkm8KPVy4qsPjDrkeBlkT74gjIYcgQBDT/srPz
tntphxQBdo0/hm4UsQFLBdr7rSSDz4lx0aguFR6FzeNWYNzx+prmWuMr4aRsZNsP
qa8Qo0hEH1RQW4EMA71HE7tz9fLXjuew+szPwUB62FcsVz+jQWiInx6PmINWhdTn
sY84PnD40ZnbnH3h+6rKMRaFag9k7JVzhXfKSGmUOdI0vmpPr931Z1xuSgpentER
8SUNaOkuzJUA7uJJq0albgP/S5r9nqCsvXZKwWFJ/Dl8SdYGncL881K/1TiJmi6l
AGBGcE/52sRx4qzHaAN/TGD65ogK1M7Y2V2B2av8R4JilMlUMmEgQJLRVOcvsr+v
HIYuJadbr6jL27rp/oyqRcA90dcrDS0qKOwBZ/XfxcYGXLQ6F3B28iMfrCQtVPSi
1X8KlqWK/H1cJRSIiJr/Yo61aP3GTYzawSeIFSiCKOlXByaRCeC33vCN7Y7FI8wZ
4CQGeMw/hMB8qul1p8mOfi8+hG9KVB299npu7tQ3Y+5PC1VwmidHzX7Wa7ZCi2e9
OyNn89sN9vFqtPxTWnVlsBZSTjj5shXvcLXfg5s9ckgr8vlgvTSGZmufr5FpSLIr
r2NAiGxhOeaBs9REx3NKcgwvddVE3DRuvKj7G8duay2iZ6Bz2ycDV6QHD4x/B3Cj
gDV3//Z3jIC+pyuzFURTREnM7PccRpVnkBWUwZWlbIgrt+IVYUODMqACUaaGho5s
AOV/6HtLAknwTtlew4ajgU26x3r/fRtOXz5lgA1rTqQBmUDyLIAuAprZjc8K9KTI
sVQV9nsKEFICabeZ0z999S02R38zBpARlr3OwdmAiGhJpW4TSF1mXTtDH/lEhkUf
rayaPovoXr2rVAO/pLmkozfAybWDvdgwOzllH47AKocNzQEsNlLYfmdV/rBRYnw5
L1/yexgtQ0h0bTDpkEfmi/7432QTAQM3wFLy28BhClFM3/Tgf1jaGMRKwldUzvrq
NddNk4b3tW3BAUTkezHgfKQxhLVYzZEeqNolXLQc2+hL3y6m6qAXgS4Xpob7IeuX
8P1WikEaJeq7XrUALuUDnXIGM0WvMm48agB6aoySnGytzOoA0IwDDN63Lr1gRqt+
xi5OK8VwQyFuKx35loG1zAAcUWWl8GNu8xz1XW8D/PNFV3u39FoxyuFLRxIFZV7t
GixwYOCzqXKL9rO+l9JwS93pBQA0pGM4i7hnaM7xibHz9VpnQGldL0YouX2UJyk1
T6Z/My0IaCeT+WObaji/UFU8QZp9EGgFJKBLkGvrpfqoYCfaAfFaW00ATghJAcg9
j4dZBxm1ZFF0NI6OI30uq4MLRTyC7WFYxRb6Tnjz5yB/tNWwGxpKuf0nODA0NnGh
AMqMiIKP/O1tukthj5Y9CXYtXchgISPU0021XhIWZESzPz0ObeJtA08FfbwVYtSB
ifzGG2cvImFR2M3owUN81dxg5P2B8SWbbZGSeIe3/lMM1J56iCBt1gqkZWvog9T/
CMWGDW6GC168e9Fv8ElNRw11jh1WTc87Ik85xA+IDrrlPmTWtErp/gUt4oWhGgG8
eBOlm3bKDPsliV9vDBt34sKuSJFgIbu3Lrjhj78xem/LOUc4B6v3g/yFO6SoUUAG
9efx2Ai9nieEAgB2M/ILMcZuz9d9IGVHgF71zXPhtuhmogu7ivznRWdwdviTwti2
39xAn2ra8b0R+Nm4//YgUH4VyY3E8LVrumqs76G2BBQoopePmsA8sl0P9hRwcgY6
hsBTPQJFKsgG45+m+Doi/9yOcGrxDjsOUbo2v+NGXFP22Y55LA6IqiaGfYchwgxk
eEkDork31xZcEjj/pLaxJcu59sd7LublL4f6RAJ6XfoGdgCc9xPE7dXf3huhBYss
2MIDN0OJSkwStFWjQBqJIQwtwKIincvrySyKD7Bs8/yHJgzMyAvRDFihu0O2gcyT
/2KxuNgvuTWUR1zD23Nc4/en5TB3BLkghM0zG728orVZ2bIRsZ1Kj8ZJWY/EJd9X
Aix5E8s8Z83oPp8DT/T2//YHPPxIpPTS4H3V07sdAjIu7O03ZpDpaelwQ1Eo+GZY
D7nC+ttlJTK92ZDgqlbCph7r+UNrCO8vvh6KJVWHWgXaD3XPtWcJ1JGzSsm9OD7D
nIREKu+djRjEGoMiC+ISlal214J4HalZuEX7Fh9vmDnOUvBs1GSte6UwctQV+sx6
00MPf8075rnZvFPY5Oft1UkmNRM/fi5AxtME5U8QeImOYirr55pZ2SA6k3ZDbeAv
6kzqPAkpKoufPR9MVLP94nx2HXw0blv+Rf5hP/KvTUj78if4CJJ/nPF2mR9KWA96
jthR5jBhZnahEYTHs7Q5d3CkVO7gbfo/n2MtAAFV6txjMbb/S7Fyl73sTFpwCVAZ
HchJK6HGh1q00RamDxqSW5I8ldO+lfwn4OoW+eO4kkvXgx49B1afJbtSiBuW7+Oi
1eKx7ci4LzgdQZCwFDmDX9Nbb/RiB6c/zRi6GC8WrXR70uqtxtr9F7K9IrQwRY/4
CF9TYuosBFm+xpHJGrmMtT8cHDWj8gCrC8vYWBWlo08T41UZZk8s9He5nkmPIj/v
s9V51Y6FFmZMCWwARcp0AL36biGrciy0wtwP/pA3arExPORrU9pL51zLRHpzg2Oy
yjGUR1vtcEhc9HET9Zuty5tc35zPtw+9XQ+IdHwJ8kkkjU5J0DajI0/AnnWRt+q8
ORCkpGw90+nGntlbAk/y5N7RbHtoTvxSHImxuPk2LpXXWkxC+tYBbEJcNSIy+OIq
yznyEZFqhSNExOManQO4tIAYrC0y05bgJzZTdg8bs4VNQJ3nSvAsAL1nEsGpCDcK
cP2LjK2hGZrswbe2vgY+GtqfGO/aHaLJSaTuv5hqj7dn5QAcVvit6ku5Fo8w/9hn
5nDN8FcdDcrAwXXU5L0vd5a0YVWmQuJUSCdWzC9EfYU224na87JbN3FHTp0OMDYO
pj0GDTF56P5ryZWCaq6Bvi1jgq42DSbFnQ27/SueDGkdtY6VzHygff8jOT9F51Qz
k6SSr/DtmyVIiGLq8pAn2ffQWb4gnxyccnutlKpIA0fqHlGNb6WMqIY+IU76qnLv
/xq9h7Q5K9gIJhInyZoElJDhdm4CAztuwsqlnnLtLClcRtUCzNAqo0unn412/hjG
8w95loGHmId5sLsN7Rlu3pjP1MJNDNNMSw/N/KxCqgYcsVzIp+viTSXtMjKNETAA
sXwnPbUCO8cfocdJCs+iqbhFlGg7YnXMCFgXRs650aglRjv+vsieEOgTdkzyyqry
1Gh4SFj9lR2v/Hu//iPenWMu03wsXQAxxB28PTv8l5pkBPc55iP9yFnO6CzuhsFa
x4lfwusLeGlgVhZFNgYyEMMsx4emynYGXYsmW446b7fBVE7tXqpi79Vz1fjYiv/j
qXaNJPFaxV7tb9tk/ZfXv0OeMuDJvjhI/FlNx2C80T+fLnJsxlXaoorKM/+DmXpM
0npvrbD7VN/7Efo2qwLJjJE9JfSvqzw6/Vh7sYk7/8ZKlIfTn6gkBrpv4/psirQf
HDWP3fIDdfjAnBQI3wv5xmezlJ8ZCKTkbHpypbzhSsbnFUQaxV5FUY5rECTDWaqH
8z4YLe+bgNAKEw7WogrDr5VB8+enpu5n7eDSu7BqjVb3aqthWySqEQMyVVbaBUFj
7bC0xNvaC23K9i1AaCDWhmpKnP3plgPJq4PtMPxkRpmmHBceXCx9Yx3iyLbNRJJY
kgNb1k59NaKBZnRLFSHN1Qj4AbfgC/T4HeFk36gC6XvioW5YRtbTYl5v5d2FhDHA
SCi5Kr0NEsbZ5xf0g8gQtaXBpQnZjkh2WrjuieGwH62qIvSMgHK6YVTF67P1EBbq
RM5ug7vSsNGKUO1fWxKwE9A9dXPY+mztn21ecyz40zIhmie4MrafAV0pXu9UnIyp
TvbN+s/Z5m8YY1ptBCYywrchIXto1qWj50WpDp5ONiKOTVSNnxeqRke+srStdcpi
ToE3jP+8RuvDSIpTry1ujvcbt+FrTIizzLW5jKgikBmQCTyb+COJ5zg7a2lQ+jwJ
WYTkRJXcoS4xtyMzFp95rFZqmWpejeWDWUTGqxd8lLyfG0ijHV/d82jLNcjtpdv0
KnqxiREeJiB95+P3+miXB+ZCH0Xjl7/4ITk9ZlYYEDTFqzUD0jGWk1eEKzOXf3Sz
UFbJ+fFGtXh/yrGpoABo85x09sV4P3U+3HmDwf7eDuV01z9eA9/pMLUKZg0w4mNS
xFkYLDyiW0WlegaauErT0+HCLhKBSbJ9IbYPBKkO4ZbLTeBBVgoaYGXh5cby2BnG
if0OfGdmsiMM0IjgTgvsv08KbUgAJ1EmmKbu4/g1H13zLVW93U9A11ypAIQ0mxat
nDsIsIp22cHwxHx5IPRLe0QQNFqZpfbSW+aQAkdT6wnNin0wbKXXQ2+miOU89rzj
vxqGVoKCkwiL0Inu+fuzTthD/KL8E4MQvb0Yh8o4Ig2ojCmgN/JPbZ8QE4+wFIT4
DNR6yLDS4Gy20wQU9NoinHO6S7aPt57bacykqgxeOxDgzmzxrYIrYDJWan/cWpkK
FnXmlWdk4646ChpuhT2DU/5PjQ+JsDXjNo0vpKfjXNBGYsdbU2LE+SyVnoGyAS18
tlXny0pvQTlRsxRtdNq4y279WSQIlhYjTLwB/O/5dXRsSnjg7Q+hDkWc0XXGE4Y4
Vi4RxJqwdhpm6asALmreZp+v9qwln7mJ5M3WBM2NO38dGwmoZE362bUWDQn14zHk
nzUtnJzNVpr3bI4Yl73eEo00j9ZXZlZ/qQpvbdV+RI9XQz4gB99pclHlFyotJeOR
PwWIpoa2WqKauXXFGxqqscDTt+d/kJRDADMhggwvCbY5Ly0FoN6pv/jS7aei0V0r
p+FKQZHFppAdMl2KabViMs6CV0L+4ZgC/xfS5CzFpsl2cuEECP4ij+YB8AOprLnn
Q+VPM94loTqPrlkRnfGnjTjiOdX5eoWSWHlEYKbwgZzSWt0MsRpQoIdtnHti2BEJ
LE2FGfud66UxA9AgT0j34YCMIm6DLajK3bXOFujHkkZMV5Vwodp7aW9EGqYWHEec
uMQa7aUCe8ZtVKCHzNot1WSsL87O9Xag/gnJaJH4R7upX1C8rEyyzaqKsuK4rSmB
DuF7i7TQymevZTgGtNGKwy4eDxma+jny59xcZKAabPPAdYQOj2Ycev0sptEOMEfY
S07qVR6wULpgOkolB3ETIblF0bQSHZd+/bTlhuubHXrsrQJVSWRms/krEw/luSJA
80N5hmXjWycEXuVCvYBN2BSgjIt7CUFT5AmGLKaf1wwmMLTn4sXVhcGeklDAMTTu
W7ReyBg929D7tkEI9JmUQREOigtXmOantork+hFHzzdr1IRpjYF730DQBjoZMcjH
Thy43qcfzSBBbQtKKH1sjY28gSLVU8qljgK0ZZJhzqXXUTC81jmomdVMRf0Zpyjv
J7D6sR5x0bgA7pLrWpkihIMXP60rFdU1UxLVl1jhXnWlKj2mdeuuJaApH2/QUEn0
ZOmoa7KyYO64QHn44+PpW1L1/E+RQaUnHAC1qdZPNY2hgMzMH0skTiMXG7gccuya
3BOmjITsTIV/iTN7JiPvBDvUJbHQkP2G6HgecbQts7DAqa9bbCOOX0J0HEa9yi/W
xY/Rf3ZzHO97xguI92cS7H7w+ZAIyNTda9CEMC9aTlqfgpsG8NS03S9b/e8whqhY
lsJM8ugU8kKAd62SmEHHeNPfpitxMwHhkSqgEyLAnxYyyk7K2OSlMPYbOe87V6WN
cUiNUoNkCkRgGS12OBwxE1YwKl3Pa7ZHUWefjk787UZ/Ib2PDD+6Ip/GTJ2zlAlh
cN4NChfsyY5xQq7jGmZsxMQ2rkcnxSclS8fjiMQquAwCZLnuYlEWEZgkJu2mXq3H
ukQsC5KMg/MNmywfAuKUNk/7FDMLHuDjGfZtbvzv3HC5O7q4zQfwlGLMk05N4cKt
a5robWVXAYU/QQKRpyFni3JuSWTPWlerepUcCrngt6bMcHPgeM/0G1lE3Bl9tAbN
QS7l+2tFIoR3KJkZupxpblsNGlgj8k6a2dp1GGDO1EjHL2rEizBd0wEDw8qbr1Gi
FP1ps1rlip5imi3hhVjT3IGVn7SOR6O8SukVkEfW0m7o93ac4UZOIH/PuNunegdZ
gPg3MJr8CDchf6On/D0cq+YSzYPRiGUfBB6pXNrHGrcdF2uUpTmyeVjBP7ePIMXy
QA+Bwt9ffIbOGmQifQjyOhcUBmm04u/dhpHWhaqfp3FM1chjpG0fcTHWCNDJRVsm
QAzMXzq7MbHi+gq80t4tHO3rPtT3reViDH7VtHBRW4rcAv65pS/pKloNzgWyuZiS
Qqq2Sd9f3KNBylKKxtkkoW33BYnea14q3gSIGXpCezhkVVPYKjot3dypKTSjWFDz
PRrp+lvdqY7jNKw9OMlEw2qZx/mlx+XsMIjpnWkQDF4l/hngNf6eCwlV36YweCen
LxslE7N6eFBW4H+cHUCfmmpIZtXnIGdcwfxmdKCI6yJQqFe9Rs2Cjc2sqfnYSg4z
4OluVh3247DTGMZEXJhFkw/68ZkWI8V6X+E65LULK8Ajpzc/nwMTrIb4gznXWFOq
qB0e/x/k6v4L1gaCH5eqSmvTcfo2CvUZb1DGIdzJ6Y44yNOwGKFruc9u6m/cvrgp
S/wUQFpUQokJo0Dlrb594/bnSNeDi/78Q+gwB3Nmr8G/jPphsMKPdGo0Gu9z2/Cu
3END3ul+MCSvZXbGAb9kyuEi/TgRi9KNpXCja8MVFt5qNL19AuXhLQbUJfGxdt7C
UIE4nhDNSEDZRegkkDwnLdfnkiK/BpWwvylvL1/cy8TLPXq2ww0B6MFlG4AfZXb0
MbjsdZdHwC08Qumtjwjwqyz5DZdBqPL+kxp6UT1j62b4meNjcHcsZfpm2Me6zUyH
wTn7T9Ol8iCsDeCbhBsqdSt410HcsxlMLT25NpSAX1GyxRJrTaQZPgLsZe8uj/rf
G4wfa7khS2QT6dmhc3wsnYoenCZS3f0Ic+oIQVCp00orzu1LUkNQV/R25NxQr805
PWrMkNNWYnQDD0B0oyy3uOgUVff09fnMklhZkTpcx0yWTADw6HxoGoF0WbcB7R3v
COa5BDV9tNCCD4MTSstFIxSq+tBXWKIh5O6yTi3jyU/UxTa1rrEWzDy7jrlgflAb
nh948xMcr1xNXUaEHNGvxAc0hlWt2DGJPViCO3iK3Qz64fczvLJFiFBRHWoZRuLk
ywasl8dyDxoN5+yqSA670aE1Vu75vvQgS1RvYkekVS89umj6a6Zx5CHIHZiXvz+w
7P8Kj/GWJtdQtlvoNtBUJ0lwPHll3B6DU+g0JpJs4729lzHvXQDtwN2h7qHI+BCV
lFIvi+cPtz+JPYLtZ6JctKzcRfSjoA9ka4zrqKy/N9tcX8+YogmF7ZjvtueDGQc2
eCcc8hECoNN9M7E5ak6QepZRLU9YeswPwyZ+dUoCc1u0y4FLhOR7UzfuVWXKZRkh
3GVizOyEIN9RqY0kUebFOKW2DXpovs5c9U7gnpdcwuD9K26Y+7OFBVBYIz5exKFC
zTl0xgH+jfhpCjZdf1lV7Qh1UzE//6iuMrUkgwSlKVVGmfiHbhQpC5If927t6tte
/P+PSUVwHwZibL8sGgBDcp4n2+4UYKJJXQwhlvuoHekIUjCu35TeBBTmFHBDBYnv
M40XQJOGx0Jym5eNLDVe+0nuAZVenjHsolb65rooMhEI3Ehv4w3h0rtr86+HFO1t
mlOmRu7kwfQhmBoPIDOGoqCfBLYi12qFCRf1Dj9CjWT0IzKkHJF7IyY4rwjqCKKm
6LAARS0oGhgJYRL82yIvJrSwVVGrAQc+kI0yIIiUwdLbyJcCXq4938uNUr4L2hsi
Gr05gSwWKVqkGNgSPT6hP8Fy4oYMvTAEn9KgkU8qmj7t6Tb1Q2Q3uplG4ly01N/U
K/kGoZlUiotG19BSO4qmy26GhWqeldWqgjuWeJvtViokPVPCiewD6XZola3fDiov
rIJw/oaO3AvTPDan8B07dks4K500UTDOhPklJZW1VKz+GloYq6aQx1hzeigJos3k
VoBMLv8g2ep0C0n96VwY/urGiermTWi/ea42RIOZvwBysk0VtYjptwug4nv0bBT0
esauDUG0lNv2rXnpzQx/rOWM62fPohlQZCelyX9dX61V5du3gtuj4KfVkBJhg4Wh
QeHd+Bcw2eGIk3OFYtfNbRNVrJLMqzmKyE82TFdxyFD1ZHcrrTlBbUWsUfR+JXbq
6xNuBgnpFxW3LQBNDOWefaJz7B8qz+dgqw2mtmlzJdxDBaY2vV2WSao896CjQLus
CfU4od/p+ZOIiCi34Q6S51ZW+P+HccMWbtfYQ9bl9Pj7aikBxsaseO1UrH9uh3ZK
rvQaeq04rpn1RNP5ass9lQf0kxhtZNBFbtawndJLVEZN7fQUa5Mk2tS0lbt8IKeo
sq7HDFF0TlGZO5cumP8vxix5uV9AmIvi+btbVgUkMZs=
`pragma protect end_protected 