
`timescale 1ps / 1ps



`define FRAME_TYP [8*75+75+75+8*4+4+4+8*4+4+4+1:1]
//------------------------------------------------------------------------------
//本模块是演示测试平台
//------------------------------------------------------------------------------

module udp_transmit_test_tb;

//----------------------------------------------------------------------------
// 全局复位模块
//----------------------------------------------------------------------------
glbl glbl();
PH1_PHY_GSR  PH1_PHY_GSR(); 

//----------------------------------------------------------------------------
// UDP帧数据准备
//----------------------------------------------------------------------------

   frame_typ frame0(); //pc icmp
   frame_typ frame1(); //pc arp request
   frame_typ frame2(); //pc arp reply1
   frame_typ frame3(); //pc udp  

   frame_typ rx_stimulus_working_frame();
   frame_typ tx_monitor_working_frame();

//----------------------------------------------------------------------------
// 测试信号和常数
//----------------------------------------------------------------------------

// Delay to provide setup and hold timing at the GMII/RGMII.
parameter dly = 2000;  // 2000 ps

reg  tx_monitor_finished_1G;
reg  management_config_finished;
// 被测试模块接口信号
reg        			key1;//全局同步reset
reg          		key2;//部分模块复位
reg [1:0]TRI_speed;
reg                 clk_25;//25Mhz时钟 //PH1 25Mhz时钟 EG4 50Mhz时钟
wire         	 	phy1_rgmii_rx_clk;
reg         	 	phy1_rgmii_rx_clk_125;
reg         	 	phy1_rgmii_rx_clk_25;
reg         	 	phy1_rgmii_rx_clk_2p5;

wire         		phy1_rgmii_rx_ctl;
wire [3:0]     		phy1_rgmii_rx_data;

wire         		phy1_rgmii_tx_clk;
wire         		phy1_rgmii_tx_ctl;
wire [3:0]   		phy1_rgmii_tx_data;
wire         		phy_reset;

//测试模块内部接口信号
wire        		rgmii_txc;
wire        		rgmii_tx_ctl;
wire [3:0]  		rgmii_txd;

wire        		rgmii_rxc;
reg         		rgmii_rx_ctl;
reg  [3:0]  		rgmii_rxd;
	
wire         		phy1_rgmii_dly_rxc;
assign #2000 		phy1_rgmii_dly_rxc 	= rgmii_rxc;
assign 				rgmii_rxc 			= phy1_rgmii_rx_clk;

assign 				phy1_rgmii_rx_ctl  	= rgmii_rx_ctl;
assign 				phy1_rgmii_rx_data 	= rgmii_rxd;

assign				rgmii_txc			= phy1_rgmii_tx_clk ;
assign              rgmii_tx_ctl		= phy1_rgmii_tx_ctl ;
assign              rgmii_txd			= phy1_rgmii_tx_data;

assign 				phy1_rgmii_rx_clk   = (TRI_speed == 2'b10) ? phy1_rgmii_rx_clk_125:
										  (TRI_speed == 2'b01) ? phy1_rgmii_rx_clk_25:phy1_rgmii_rx_clk_2p5;

//----------------------------------------------------------------------------
// 被测模块
//----------------------------------------------------------------------------
udp_transmit_test_sim u_udp_test(
	//时钟与复位
	.key1				(key1				),//全局同步reset
	.key2				(key2				),//部分模块复位
	.clk_25				(clk_25				),//25Mhz时钟
	.TRI_speed  		(TRI_speed  		),
	//rx_phy_interface
	.phy1_rgmii_rx_clk	(phy1_rgmii_dly_rxc	),
	.phy1_rgmii_rx_ctl	(phy1_rgmii_rx_ctl	),
	.phy1_rgmii_rx_data	(phy1_rgmii_rx_data	),
	//tx_phy_interface
	.phy1_rgmii_tx_clk	(phy1_rgmii_tx_clk	),
	.phy1_rgmii_tx_ctl	(phy1_rgmii_tx_ctl	),
	.phy1_rgmii_tx_data	(phy1_rgmii_tx_data	),
	//phy_reset
	.phy_reset			(phy_reset			)
);

//---------------------------------------------------------------------------
//如果仿真在500us之后仍在进行，则说明出现了问题
//---------------------------------------------------------------------------
initial
begin
	#500000000;
	#500000000;
	#500000000;
	$display("** ERROR: Simulation Running Forever");
	$stop;
end

//----------------------------------------------------------------------------
// 时钟驱动
//----------------------------------------------------------------------------

//phy1_rgmii_rx_clk = 125 MHz
initial
begin
	phy1_rgmii_rx_clk_125 <= 1'b0;
	#80000;
	forever
	begin
	  phy1_rgmii_rx_clk_125 <= 1'b0;
	  #4000;
	  phy1_rgmii_rx_clk_125 <= 1'b1;
	  #4000;
	end
end

//phy1_rgmii_rx_clk = 125 MHz
initial
begin
	phy1_rgmii_rx_clk_25 <= 1'b0;
	#80000;
	forever
	begin
	  phy1_rgmii_rx_clk_25 <= 1'b0;
	  #20000;
	  phy1_rgmii_rx_clk_25 <= 1'b1;
	  #20000;
	end
end

//phy1_rgmii_rx_clk = 2.5 MHz
initial
begin
	phy1_rgmii_rx_clk_2p5 <= 1'b0;
	#80000;
	forever
	begin
	  phy1_rgmii_rx_clk_2p5 <= 1'b0;
	  #200000;
	  phy1_rgmii_rx_clk_2p5 <= 1'b1;
	  #200000;
	end
end

//PH1 25Mhz时钟 EG4 50Mhz时钟
// clk_25 = 25 MHz
initial
begin
	clk_25 <= 1'b0;
	#10000;
	forever
	begin
	  clk_25 <= 1'b0;
	  #20000;
	  clk_25 <= 1'b1;
	  #20000;
	end
end

// clk_25 = 50 MHz
// initial
// begin
	// clk_25 <= 1'b0;
	// #10000;
	// forever
	// begin
	  // clk_25 <= 1'b0;
	  // #10000;
	  // clk_25 <= 1'b1;
	  // #10000;
	// end
// end




//----------------------------------------------------------------------------
// 复位 udp
//----------------------------------------------------------------------------
task mac_reset;
begin
	$display("** Note: Resetting core...");
	key2 <= 1'b0;
	key1 <= 1'b0;
	#400000
	key2 <= 1'b0;
	key1 <= 1'b1;
	#1000000

	#100000

	$display("** Note: Timing checks are valid");
end
endtask // udp_reset;

task udp_tpg_reset;
begin
	$display("** Note: udp_tpg_reset core...");
	key2 <= 1'b0;
	#400000
	key2 <= 1'b1;
	#100000
	$display("** Note: udp_tpg_reset checks are valid");
end
endtask // udp_reset;

//----------------------------------------------------------------------------
// 发送UDP帧数据
//----------------------------------------------------------------------------

initial
begin : p_rx_stimulus

	// Initialise stimulus
	rgmii_rxd      	= 4'h0;
	rgmii_rx_ctl   	= 1'b0;

	// Wait for the Management MDIO transaction to finish.
	while (management_config_finished !== 1)
	// wait for the internal resets to settle before staring to send traffic
	#800000;
TRI_speed=2'b10;

	while (phy_reset !== 1)
	#800000;
	$display("Rx Stimulus: sending 4 frames at 1G ... ");

	// send_frame_1g(frame0.tobits(0));
	#800000;
	// send_frame_1g(frame1.tobits(1)); //pc arp request
	

TRI_speed=2'b10;
	#8000000;	
	send_frame_1g(frame1.tobits(1)); //pc arp request
	#800000;		
	send_frame_1g(frame3.tobits(3));//pc udp 
	#8000000;	
	send_frame_1g(frame0.tobits(0));//pc ping icmp	
	#800000;	
	send_frame_1g(frame0.tobits(0));//pc ping icmp		
	#800000;	
	send_frame_1g(frame0.tobits(0));//pc ping icmp		
	#800000;	
	send_frame_1g(frame0.tobits(0));//pc ping icmp	
	#8000000;
	send_frame_1g(frame1.tobits(1));//pc arp request
	#800000;
	send_frame_1g(frame3.tobits(3));//pc udp 	
	#800000;
	send_frame_1g(frame3.tobits(3));//pc udp 
	#800000;
	send_frame_1g(frame3.tobits(3));//pc udp 
	#8000000;
	
	#8000000;
	
	
	
TRI_speed=2'b01;
	#8000000;
	send_frame_10_100m(frame1.tobits(1)); //pc arp request
	#800000;		
	send_frame_10_100m(frame3.tobits(3));//pc udp 
	#8000000;	
	send_frame_10_100m(frame0.tobits(0));//pc ping icmp	
	#800000;	
	send_frame_10_100m(frame0.tobits(0));//pc ping icmp		
	#800000;	
	send_frame_10_100m(frame0.tobits(0));//pc ping icmp		
	#800000;	
	send_frame_10_100m(frame0.tobits(0));//pc ping icmp	
	#8000000;
	send_frame_10_100m(frame1.tobits(1));//pc arp request
	#80000;
	send_frame_10_100m(frame3.tobits(3));//pc udp 	
	#80000;
	send_frame_10_100m(frame3.tobits(3));//pc udp 
	#80000;
	send_frame_10_100m(frame3.tobits(3));//pc udp 
	#80000;	
	#8000000;
	#8000000;
	#8000000;
	#8000000;
	#8000000;
TRI_speed=2'b00;



	#8000000;
	send_frame_10_100m(frame1.tobits(1)); //pc arp request
	#800000;		
	send_frame_10_100m(frame3.tobits(3));//pc udp 
	#8000000;	
	send_frame_10_100m(frame0.tobits(0));//pc ping icmp	
	#8000000;	
	send_frame_10_100m(frame0.tobits(0));//pc ping icmp		
	#8000000;	
	send_frame_10_100m(frame0.tobits(0));//pc ping icmp		
	#8000000;	
	send_frame_10_100m(frame0.tobits(0));//pc ping icmp	
	#8000000;
	send_frame_10_100m(frame1.tobits(1));//pc arp request
	#8000000;
	send_frame_10_100m(frame3.tobits(3));//pc udp 	
	#8000000;
	send_frame_10_100m(frame3.tobits(3));//pc udp 
	#8000000;
	send_frame_10_100m(frame3.tobits(3));//pc udp 
	#8000000;
	#8000000;
	#80000;	

	wait (tx_monitor_finished_1G == 1);
	#100000;

end // p_rx_stimulus  


initial
begin : p_management

	// reset the core
	$display("----------------------------reset--on-------------------....");
	mac_reset;
	$display("----------------------------reset--off------------------....");

	management_config_finished = 1;

	//------------------------------------------------------------------
	// The stimulus process will now send 4 frames at 1Gb/s.
	//------------------------------------------------------------------

	// Wait for 1G monitor process to complete.
	wait (tx_monitor_finished_1G == 1);
	management_config_finished = 0;

	// Our work here is done
	$display("*********************************************************** Success: Simulation Stopped****************************************");
	$stop;

end // p_management

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Anlogic"
`pragma protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "CDS_RSA_KEY_VER_1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
Xl3k5NpexXK+Rn2vC+7vnXTKVhAWnoDFKVqb2OLP8/AKdqtvNbOHT7lHWugEMYZ/
mLGBxji5Orl8AvnrzknvmlajZyx+D7cZS7FRbdJaVUfeLRXG5fbE4Lo7YH26gtdH
uZilXa7rCDeFj171DzAY6CnDgMmPvVAFowhNFo/Q0W9I0OydDaF4Pi0bLiSSBBhU
jGJ14ttDrOxnh0NOPZsgWFlqAMgye+otdXMFOxaQuTTXUmKTlS9A0ewcXzRdzQmc
nNmyh8cUyKJc4xdDs8wpIO9BYOB/zriXX1k1/e8OZbRc/iORzf2LH+8R9Kv80ZHs
OUwmk11bp673nJsqL48USw==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
IDrRGmy7j0t3shucCpcC7BAMZXkM8mX+oB19MHs2bsaZVPfRSMDjjYsTTdOzt2ZZ
0ISbw2El2PjTwKqFHIUHofDeEY8dK9eg4fWh1RGBzAMi/MJUoozzC+KWkeQwPMCT
MUcp3uBUB2trklpghFNEOvTgn3sTIYVFuCPvKgWfqhg=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
DpLeC60oCmK6e0HXnRVnNjBlYKXtXMBIB+Jouf3YzsDF7dpO9vgzVsGWZCeXnFgF
BAzGCS1y38t6SmyuYfM1Dhwit5KaqxXGq+IWLqbU/uNKKTolcfXYlVBu17enGXVt
e/y5f/hnkdhm/6eMGSQqQfU9rwEN6YxdkvWkwKV7l7sTNtRaCSLOPrGUM6/2tIiw
j6hseRPjwZ1gHcEutIgc/8aV16dYWVkwNif2Ta5lq7wiQxynii/a2JN9cmgGQXGu
fLk7NBLmMUNBGBkKm8lOD2y3Yl8oOS6djtYNDiQyUCr2GPSUqGIrvj72jvlYfukF
4D6zt/1zIj6/BK6GBoMllw==
`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
mg/EWBN/YbGSh5U8C2uySUEF5VBX9CIAzuCcULXEbmOX5Hb07yMtg500S5Un9ih4
yWdspLQgBS6g52ZU+1DnPCA+SagGlzgSn2kURvfBUeICmWHnbfsDdFglRbk7yo4C
WdqGKqpVz93zHeGBWKS0dagbbANhfCHRuhyCg0/BMvE=
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 36448)
`pragma protect data_block
cEkxdnBlTzM3Y243SzV4ZIPDqZ51L5aPcjZGmKBe55XejdR2PqgO0fTNG9nYyn+O
bKuHzUkMZyfnz2rTn0ftJGBWAzDOxsPMmCcvDGhQncIzg2lLshUsNHtV/otcNsfA
4cTuy0pjsQvxchxk+YZeMXSw1T+wNAU8iX1olmZCC0/uLSZSoNDF046rty+ErKL2
rvc8+/BvZiwRUU+hXUDtYRNFddJ/QeQClZsyhuiF/XWgvGlurCn3EsqSOl9o2m79
7kRkjYwiYER1fKIrVgne/45qx+J7BX1pB7BV6BeMz/KlkaEcYbq1QRoGh0eU461V
JGabift6hE3zLitgjUyjSZG9CNryMWjdy3KJ7bZLtg5DcZYDet6KjaeSf81lEPEd
y5mD184BVvosqj4ZHaHv5kH2IUKEV0Xw0FMubKGyUu0JKuWeZ31+hEtoIuAiH50o
YWpmKN/Yg/iqBS74/gkCxH0C8ye4y6JB6RoEuIxfyRoajhjSOG3+7WsyiUKZ/trf
5AxEbXunoOg/X4WJHewwtwaMAnWic6daXh5s4GnsukN15lf4wXZG+MTcCy5fsRvZ
ThFLmCCbW73G/KgHUlWGmCHNxGR1bWLytKgki56xaYmWXoV7ts4vrEVnsfPhEn7x
llmE3k3Dx3QUomrpA+x0ZQllZ2M+u7iSietNTJvGF+6hB7eYYtxYvIT5FTxGM4um
hJZ3sPM5ee4C8zK4EfBiTnAOLj9TnRNPCceEFZf3Nzut7QXey0t8udAyIG3KcUXO
dK5npqrrWk7Lh6KSa1ZSVf9zjApWLjkbagm0mXj+z4VYeYUqdnZDM2pYutNXk0GO
bEpj3oFhalFBWKzBYV9tf8v4AHeY68ZZaywlZodZPOXYR8JWGWR0yePSFxMJwLNj
2BkP+j96fLGCGTl8su9uADwKYhBF6oALrerKOhZF7PAQFyc5hqnVlHuHQEtUoHXF
D6bFQvEBO5nEsKpHgaeNkjV+aC8Vw60YdgedhifIuAI8QAgAEpI+LNgupc/cbBIA
mm+Sric6gIPnH12VRbfoITKrFV0wgYeniTkp77/WOxPzoELF941+tP/QKtwZl6lE
jCTTr1ucTKhrxfZRdsxJv6Y7RVVCpu3aM3QULlSOYlt5h9v5kZao4XI/0NSBVMW4
koaf/C/cKMejNjapveviiZTCRmuavD4x2TkBByVQOh4JhcbfblRHctKZo98MoHJJ
k3C/3SpgcxaML2w598TtNV7T6GVShDYVe3iewM3DwvkLoTVto9ZWA/kaofOqGN/B
6HcAndUa1FUkfR+8um/iXcOG0XVd1X+WAIkpsd/KGZEOmxX5S4GpryZRKVGE9dAi
1Bf3LvDztZzig3ECwegF4oXYAxUGWemnn1CN+p/HXqYf8w1tI7+GN1CWpg+JTkdy
76UlZ8WvfmB6JCeow3ZSkx2ZN+EFlh3JyyViuWAMb886u5zp2YB+/Hua8G4L72F2
PYNQBVKPZrztFiwFvghct7i57e+E+2kIyZ4GrOx83GBLQXIA0wYzZOYeOeijc188
HmnGffwQN/CiGVj7EVVuyVFFSrnojXf0X/fENs5cBHgc0Yq/bQrASkAf58FiJIz9
x3T55ceY8s0/Zj6NoUpOTrJ7CFAOxDtHkOVnDnI6n7zijOtDPR5PTbaRuaJGx7es
m3fPXDFeRJj4TeiJuCURhu2UdK8/NzNZMDEhOWsvFQNlk03pIwGCqDyM+VEfwpRH
laIIPJd84HcIpfQqUKUZule8w4m08q+SgusbgizliKkCMXdnt88kTov2kDel7F1t
WrSOb73VTzladKSxaOhU8YA4zzNLtTawF7dyKBT25mcGJQ/fYohMZs8kuCSs6a2O
wBAB734yp3ZZU3b9aXx/eglLPua1iC2rCAubPUGnOp2e1Bay6zHmXq5ulCJa9M+E
VA2beXx5WNkJ+UbZyTUEuE9OPUG9bEBgpNgz1RsZ9tPg+bz1oE809amOCoJs/XKg
UoG3+o4hUtSTdtK/DYBDK7TFGTtjIirHIaJ27nNxXi3PPCAY0q4FeltnVhAZG3m8
jGMjt1aiHt/NsnA8KNXfoIgOZMIMqJMl6bf1ipBOuTsmMPyIVWxRTpd32scuARX3
1ymPffESjKeiXH7SJXvrSTY7F/x7XZuuVd8SMRWLxpuwx9N2JRzj9uTu9IhtY8W/
iCQ7zxyJSo3adtMwB1ntJsq70+bWy6DsfmRfVvJoceU02rL03X8ty11ndRC+E8Cs
5S4aH7r9EvKCG/bFvn7NF828MG82e4XEeL1XYfPC4G7cEHTqOzFMkR0QwOjzPF8j
QZQAi9sPmFCdEHdlCMlwiAkZQU0puive+iPVB8hXUKaUHrlZfRhrYSGZjIp2zj/v
KKz9DHGCmpnB3+Bb+0e5oNHNDt0Bm6k4scTBfri7I5WThFFCKd0uKRp6Vn2+ERpU
oeHpvFyKeRLPpPRqmcohtMbRkUQF9P3dUlmGcM4k9M6ogWjuSyISAS12IEj39Gdm
EF+HffO58H3q4xWRZpI/9oIAHP/WK08jgjSlp0xaR69o6tvlg3y4COukacrKsFho
huc7wupWiLJh7k2f/DHpIgEtFl1/kNfRHVSGiBv4S6pwfWxHcNdwUx+uQpXj7mlB
3nmsowA69PfbygHSeZwrtdgjDnKSEK/0urVvx2DFrzsNGRNxymxtAczbVguqZlnL
m5aG9dFcGQb3OT87DLvSCAJe+GBPsPztJb4J77D2dxPGUQwKDGgbA7vI7Ob5B9tF
V+IO36YfHIa+NbO8pnKEiplXwdBa3NmFkie3U9q+gpBjqsfVoyCijsf0aw1sEYmV
XXa114TGrHZOg5g2j/qy3861zESgGKZ9yGMC77mpQtZQ+9pITDKMdSzVsOwef0cV
YOIAqrIDtt8P7ca7mRiuJsuBFY5rWyCLDVgp1eVBD26rcQYdsT+sVl8lOB47fGNI
IrCUHnxLdxNUJ9l3YWPY1HfeP1InC6uXrHZBJYgr7Pxc9D088q7pRUdWLMpbMG7L
vVbSYSoiwVGsvUGA1PUJwaXOqHInQ8wtxF7thPnCxQAsKVAYEla69N1Uhb9rumb6
loe+R3GNW6WPoq5uLTT8qbcLNagcCSzCVFes+2MMMZ0RJOctwT+F1hgOsCegYuWi
yboUj+uB9GSFBjwIyMHsx4CAoAg6OFvaSG0eONk3GPmEdmbOPRwVUAeo+55l0c+b
uAErHUrAW1sTK5+Rim+fqirXQh8sh+uMY3m54MaPhxxBm17Wo1/yUT8JJmzLs1Vs
otM8wlXbFVcrCMB+O5RbAKh7eoxM38fiwAmY9DXj8zcixtxRY6Ziqjc+mQmstqvg
GB4eDMHpdD20S1RdwY8Xba+VJb+ge9gfEI7yF6UfmNesZmfoDI7b8qlVD4M90DOq
0kfpACRQbu37llsFQ2rJn3FdASTCgOyV5PxUy0DT8R7/ELmOD6BXM/ivZNd4s4vx
d5Cmf1xWQ6Yb83p07Qe/7XkT1LRyTvKFBemXS24tG6yqlxQ00bcXRScPO/v1xhKQ
GvgfnXBKtIARvV1NU73T9wLcOH/nohTvaeiaZ/4UGyI69ns5pCCDjP2c45fO09mp
ufY8CidgLGxntmrRtcO8AFODvwLmEU63Uqr/iMtT+CuKoBdPqFspx3oCvKSclKDm
LuCdJiP581DUYcRNy+M2XdeHzNDSeQzFsIPx2M4TJMtl7LkGl6bRSklDslOtH32y
ZR6ObC4zW8MoPgqWHELpxJuA8G2Vc1YSNh9XsiI/BfMk7q/YqIY/lHRMOBKn2VGH
lX4xEZTLwiFZiY0SPJopuW38/FMsaOou1wnIbQ2plXOLxNb+2SNxWrgsMBrW19ma
F14zCPWZA9eFqoVa64lBYrNGj6CjFMhLc++RwYSMGl2AJEZ9lz5GCmw/ufBOYI3L
I+6fQvKRYN/SRUPmV8FVAn371rcqDmgzpXpKVuYf5vrNTp3h5hcnAHYnaUkEJJ+w
a2E6yEhrzp5r3KrYGzbq1TDkU3FochVufu+OSRIM6H4KYqeydklhHDIRuRJUuTNW
vfbD/JW1b4PyKr0jWMkA2tXGoI6Me+6vpR9BxA4M+y17xMndKH3KJAQlUqrBvp/g
dG+2YHur4gDRr+BavWnHyp+cqx2zADnhfFs+6WpvAyLWt6Cf7RvcAIIll95sufOV
cKUs5KYOD+W+dAO/aYrVXbe+YB3jTy6azsDHw17cJQnCxJoaweogZpjMBDdDS5SP
gLYXmrPBvSSebeBZTdKFcXe5cDp0nHfBbIaWt//ebPuixV9HKa+46J2Wjqzjoe8Z
wKdMb0LWYdiC4eh8hPOaKylBNR6r/j2VhfNJQ9JN9t3MQZs3ErFINXoRKxBK1loI
U0VQKH6eWa63GuoA/u9b+2ZWnkxSPpw6gtGr6WNR9ptvRWf4iQxLETKInXUTrV2O
wKtUEJDcNWDqKkn8a+tlrplok2dL/D4kcDYkeiPAzPbfWXz4qI97dslycJSiT2ko
2DBwM+BUP2hTG3BWpb2v6mhSQG5NGrF20Q9epW4qIjv2UgNPo4tc4GvIEttaeICC
11hD4BeOMHGsfYvSxMYaYD+1GjGjvEaSso6qPh4zXwpeGA7gDwHH7tJf0G34z7Bg
/0vSteMu6Ejdcxr0VkrIct9dhczlgcX0m4+zMFTzuuhWLRXU79nLbcakWxBxCYG9
udwGChDOIlrKXvHVRF6SArSnj1IAulRMcBpJ1qakikXAjwht3pXww4WI01iUi50j
Lbkl/1y2QIkHNHi1rpszeBsTK2JK5oaXT2ZzDFgkfjGig+aLiH2gjFiNMQCqIf5L
coX2Yu6nUbPpyPDSdJibCpv9JXf7Z24Ap0ypI9H7CzjrAJo9ThHdJGss0cJFu2XV
QPrbqzlfFjopIV7KiQ00jjGMmlgzgPrWb44eJtc/z1/yl/DnsCdVFetSM7d/LW1y
8q2Qs4nmB/7k6xp4upH0y0kR9dZOCplcD9GmvZeX4qHJu5v1k2hN/bW4e2hpcV8i
Nc0TlQi/GDb6kM0Jx6hGq3dc8PVtrKIVXTAz/82G0o9aS3BbUMV2yrukoCHH2/PG
xOO136rKJz3v8GWclR589Ts2/m6LuDQNkX9SbdVa3RdhP+r8h8o9pNWnqfxj4JzV
qFecaweHPvjrSD+tIn+8fg0238D3Vf0h84MJMISRBlpgNmJVDHeCjYwkpAvPUWNh
4nd6YPGKBKC0GuzxfU+ZwsWUhS/EmBUM5GBoEL6RnSidOyKe/olPrGl+uT6PUi2R
8NddToXtAcUolxE+wUUgsL8dCoKY+TrCsHb+nZkYqMwySPDmYLiQLIbq1j/p0Cwq
svdOYDryHidDfh3R2z021v7FtnqNE/CIFuaYyyBCp/URjb9DcSZsgGtYfntas7kq
I7nezvtFoFl1lYqesEH6zlv8UVCN4GptHdffCJLUAWX45fjEuQmMhCZatxRVAQbC
3QZEwAXNwkjpGzOGHpyc0STuF5ea131a/5EU+z1k3hxZZ66wBXX9h4ZL9PpDtRRt
X4+5W/ATalzuPXzbrvyMjR1I0xp4DKrS1Pc+er/Xb6feg9lzzWqe0/Xhm5CMh003
B4gyKeUmAGGGXoeWN932rBJHIRC9s+zyZ8KtkrTDLJ+DtqkRWUFSmbjFaPqgW3S+
r8EPxG8gCPMG06SXnbjk2xwARs+SA6GpXXDG/7fVPm9vs/qw0zYL2/vNolUNo4dy
02yC6C5GQZpOJe5rDs7MciendrCdLNxsKJupvHXhbLFAZIjqRqOUgBvBORZjPwr1
wcxq9koxFnW3EfqO93PWffzwvL7ygf8BW2fB4+hExav+XMr5VRoIqFfNdZJOaI0T
F7zyYBfURlOjlkmP0aD5e8UeNstu7/2tgKUpmKOBfLXngn7hZmCb+u8rnaWZvi+7
LuxI3qRzSGUqIyF+OKKKXaOucgJDkRz+WsDsy+eBpPMEa5/Fw2lzlIVRHl4ndeDD
2zNLcUWjqK0yIWzKXFMG5SThWaAdRT04bsI531BWRUhfN8sDCp6xUOSI6xtN2WCF
qfoGzSP9AnjQK9adPMfDabs8poU9vR66ePe84f1Sp/e2aSl/rDxOUvQNIAaHD/f5
NeWpi0fb5yB6ujWowp4wIXT+K6b+6CTuEN4nIb27ZnIRJdtFONLMOk3IIEtwUNXO
kq4O8g67siiEczeRxYHq69D9l4nNxliXtd05TPETVgxS+203KZSPG7nOOxsQS1bK
d1mEAm9rPgLwlbpSIT9tO303KrpXayDDTxLACOnNHhn/2rNMiQWGqS6AWr3Hu7o0
nFUEy+O46tEwtHkUR125JCcdu5eCHcvIzRISz9V8Qp9349wcWP198MA1DTqBXzU2
56AevODDs9B75ZVjd4iaXC+XWUS8PbzGlv4pJ+aRIJTlV9Wnh7f+AGkDcigE/iQr
hZCMUXjzjQ9pwJRhaLFFTR0TeQAyWzsW2A6i3axP+fYh7+4sHPtvNGQRFvcHERPm
FdxIp9BMeZz1naP9szEHxncowConRPmJm3chfwbTd5XdZRKx4eD9+JP2XPJQv48K
lVRHYoOoNRh9T3d7i/odjmS1y6rj/fJYZlbFMwj5+svtPY7L6Bb4wplG05beo9SF
d7EyDe8fmGA3td0lCGKkPw4jOf9BVkDJTL/YSZa2hmnu2eTE6JPTzLfibWcasgHp
Hh+5Dnv34TQ5Xun6AgxHPvJ8fVvUrtOGvi069xE63ChAHRUQynsRxJq/jCFAZAgv
e2vcayTMWO5mioysEHLSxVZtRwnQ+btlJq+s3t3IbySruBNlAVksv19ecFEo5QWn
x/eoUOXcuK1nPSMl0jL5lo8vwQrhJHLFXwNd5fc2fdYEufyZAJbn2yYEwr3QcGUk
a10y6YnuvmhWG9N2lIcMNwQgxdsSsJ20xlu0kGjlXCRHs2DgXaIyia8g6cMj1pBL
pSiUWpNYct0bY6eqCiHwdETNDwVXJhMRpQXylFYMa/mDvFn58q757yNUonUOpuAN
DbPVXrp3cRNMui4e/FVqw/29Xk2S2G3gErjUCvOXq/mb7y0ru1Q8c07LH7s0oAle
Hbcl00pW3SDxZXw61S64BHFgzw7tCUtPiS8FB63hMzj+Zfp/JiZ0dSNrEFKB0ziP
f3dTa0SXnmXpK380KKbReEp4SK6PTf64DtjNLttjjPlG3USEC6WTjqPVoi18SKdv
dVLBAYUQA6mxJ2qzyZhS2BpAwsTKBGJ9V6cBUeGAWC0dMOEh15Q1VwDK4Ur0Q58/
eCPfvVroq80DHbRRmoayZe1ipeIQFSrYP3mbNDEGW0Mi5tgLV5ojIxT8efxScOkr
YDWu7xRI0CKVkf3l2epmPOxmrHE4+D7Kabzbm8QQ0TRTwKqDNJ2cdkjF3UlZIDcE
JbCtM77voMMjZInsXtHTV2Q/8pCf9eVGgbuC8MNsl7CgC6nxZQHIktbQyNPejWtS
VGsamTuyCvgtY8IEwYfzMPZtI65BRcyPHNqQTfTHmNxejlBIlmGAYOzyK1qQoGY9
56JF2AZmwzY+LUsTCI+Gp28ZiKv+3yADoXVHEYcKsYCt5mRt666M4wcvQC1CW4to
iKVpcGwtQGNYd3Ajh1IFqKnTtn+NeXoLqZ0n/iL3/TEKahRONfSchyLl38INCi2G
6/6grnuCUAaWT2jTKjoFBqc3h/tSlISqVIPapSYOVwIUQJnr0KCdcQkLuSriJtwT
iGnpAOqGGN0P61Y4aYVXMAvueorZOJnTwxlDf6wCYzIy0Tw67nQM5LyTPyZXhcrH
XT0vHRXXw58ft9hBM80PknvLLiWYpjm5iyUpLslKzSk6NYYQBwrMYFttMwKEP8d5
LFHtvR3B85mL25ilsbNiwtukeEc534hIPa8srnH5/qo9Nc1DBXMHIwRR6wwsFqpB
IkbNmtvTJX2xyE3yMNN2YzLuEyQt74imPXIEUy43AxoIqdHYNKM2hvM01lT6je/P
t0AWQg/hwrM70JzYA0rUBU2a9Fl9JVuBLHnZGQsug9hOjnk+eB++0tCSVPNnb+mv
lcvAhewWglDLeKyEgh9BJZ6ZS40EUpf9PWUyEaAkkSBsKp/y2Bi5kt/SWhEaDNVj
EiUEBBHApLHy4y98fEgbOM0NLYHaiB6ADPJCrMRsgQIdyC7YCXXsJXFD71c4Sg+F
OQI0QQmnNQEDbBPIU7chj+Ad43xdyapgIjRzerf24VHysClBORfUJ0D3s6vn2Vlh
a7sm5eazQJ/xXdloKKXNpU+8ZbGiSCr819O325M7yS6G0u2wWOI5gVqugGuUxtbA
kb6dFVer0hWL4RjQ7tQUACoSMdyWFVdbeFq5OUVwYqgQtN2Le2gKRTziakRWiKfh
1LPvb7RX213/EcEfBOgWzavJhYSs0yyJVpfsjtBDrMcs6NlT1ZKNqFk7oUcT6ZXf
YPQZTV81XyFncNOdtRqWgEx6iIjWQ1SHmzt9qjrcNsI8NuNCU89vHc5v0hwNvLoc
E659itVzjDZFojDrlBmzbmPzZVM6DfIGMRKdwoChspZN1W4iSUdb5b4nxN2ZfF/F
RNOZOm6lLUx3jkquns34ArsPIr+pLqMiJHsoAiBgPm2gdYBo2cb0o0mq1XiVWcSB
vWHldAI//D5po6ZeMS4YpAQ7VaEwgLmzzB+w/89IiaSHTsobK+freDV0fkuWW26S
FuKPTDXi8cyZO76vbzNUCWVlkQqfuOA/prvFtB8HX9kdvQfqB78ZlLemsw4gSQ9/
Jfcr6WuY3HxhLh/6z2d+OmVtJlb234NQc5/0C49GxHdUzil9Ip5bTvebiEJ+fEm8
eWfLN4cDFxXEM/pz9JOGQyuL7r96u6lIH4JREmu1+faan0yRLdHQVFk84F7UUTqB
dmpT4945mrheiaek8QVpy3NpC6uc6dWz/j4zjJb8hcKaFVIBd5BkXPkYcV3gt9Ib
08bxIU9VtMZOkGFyYpDXvDxC/WBLTtJ48++WkCsFdb8vqgq5GD5/SV1yIIkNiQ5y
VycRe4XKiDRbRkD3CJ/k50AeujBVxk8hHj2hB9SfwNewrPTdKmzuQNnXtGtSFBRX
i4xy4cWSERIymcfdqD2wBF/6FN/L2BHgEJDydGkg/VFG6oN/6PC5BbLqCk+TOpbZ
cFPfuLlYmJU8BSsgzRTR77KTiqRnX/L52DpYABLfmnrTydim4lag2h8CfdMLJBgS
P45NTYcjeLmTynIDFVUxJdvweyHfuUsPtn+BrOP5mlLfb0fRhwDkMDbE66pHjumQ
8HPRNH1gZlJNaufBVTOpdEiDUS91LIHXPukifnSUHxZD2Ybc1hSh0XB4nf/pr/iN
CVK48tj0/b++yaD4VL6cQPDbQokXdaN5W4/VniqS2TkiEb5A+SYD7mugzlvNTFMJ
ubpr4rhf2+q0/nBnfzzYSqXdv0Xvo/zeavqPWtOdP0euJlHLNuRxAEslWPzBH7Az
BqgBcwViF1/VxrhvMSsgOmrnwchuEgpeFpdg5TCstmmR5+6pT9sdQuz5ow+T+EFO
wxmErgmpcOEBR3Y+ro4HtwV2XsD4HjodthjYX16o5pN8rGow57d3CFxXU/Ht6NgW
+5j9ORXwxRCxq7hIP0CnWy4HrNMfrZxwND7sVHM5Uk4IohmB5FWfMqgDuXuxV2Ju
tsvBDRa2gFl8p1sGKcc02eiFTNWHTp30pHkNRY8Ivvf07hyBussFq+iVjM2ph3Jj
UVLj7Yx1olimjURN90DQMGFabc4JIBJn3oaYi9HRRUjpdOnlgOr+b+XFUQBIMOjK
yUOtZ/3S10CdoQhHmfFtZfcGgQPj4JE8mhLevNreH11fsS6U+SVHxsEvDPBCJu5k
RgMYwcoNCk6AL0wGzF2BWAn0yfYB3oKcgOEIzv0Kz9BTLpln97NFjOVVs5rwqVob
6+/Cb5M6xOTr6USGDKjdjcjqZmec3Jk+c9RP8FEPBJoSY6bqIL4rCQC6qSmQ4pIB
ZXMeNyV0kKAJRMajDZQ5lFmMy0um6OTixeNE/7bbxdKQRP5CvydjXXZ2IXTdAB49
Alljico975kHGd9LRyZVNVNlUYCDW0KqQZ+fh0vNYeVGjZ2x9gmdHRTlWmJ7IwrU
VdJMeFw4Im/UQQRiMCWMgWucHaUi2p7hMclR4yn9ZGcSIh+nJ8nHKhyBlQgkB581
bqCV+CyYhDt+JRawoG1GUJvZ8hHMobHvgH2GKMNFg0+Eskw8g6Tf1PRX/YBNsDP4
Nb4XiDFeQHZ+Ira9HUrPaw3gAqCggMotcRwur3j/VkK95qBWyOttR+D1BIvjhUqs
Xz8CBPCx7O6eCkQXLcAigTsIRaj/35zePKImDRcBXfpDCjuQgtHD5DGGiBisJIpT
LYTOPw+Hm3QyOQIWnlZp2xm4kf/I6Is0yHYOSeFdJVjyrSSTA3mPl4AG19i+HWGF
VrW6dHXht9Hk+YYCvJ4XgrxjZpnjteOKwLClNBYIFDk0ynJ72pCF6yYQLS0J//8U
tVh7Rw8eY5mBwg0fU/uBqe25H5hORwiW1CR3q6jwky4+tsppQdcJoBQ5WjBUn8/D
dpE7QlmS9ixR1YGLDAUwCypSxY7iMyLhFrdjfLODd/6MbW5H0W5zcgwQdH9vLyU6
4+qptmB0IQAPmcWndVkM2bRARL+smYWIOaMiAl79d7HJAFFQZKfCX8eOXhXub/Z+
5AGxXj+vnwn6OTxEC1zQ0c5akDZGHlIPsx9o05H3ukGDmcoNCEef2UpQZLrmM91f
cYRN6Sii1BifrF5W3WSVEGqBxSYxkb0++1PKPK00QTGvHsr7wvnJgEX+XH/P7WM3
2MkJdzwA4G53O+2bobG7kI55HrQUqwK2Nqa0sjXhXdQs8f1Huuglm1FLL4x1QPgL
3cs6MtDCLpd7PfIiv3wfvIJ5E/Q1J8Qa9SoCLo/dmEB5BkPc7qEy/Rz3Kt6/fhuo
D8/iwJTrwUoUOzi3HOKsT3Geek0X5F7khVbile+QTx5BbjJUXqFll1YDF34CCFjk
hvh/oPVI4+tVALMMFjODjaiv2Z5YtXaIxH2hLfXEZCkEHZoxpx82PuQpwhEYXN4B
QMmSIN5CM80TGMlJMxU0FxISGdxWqOaOcjPrbrEdQvc52Ks6sDPqTyhbPYL7shsU
2LGyyvDfLwiIH5lCXhKX9A2MkXC+OWm1T0ttysq19sL0T6tvR7LhuPb9k7JDHR+i
0/6hyMn2R3FBPJ3iIhpouJyZN21uWbd6cPuQnYiet6txqudfatoJc39cQHsLz0ir
2fyBbQWg6Zs8QrRaOQumRZ7fOlyLBE/7kMLZrTRbtJZMGx8HJ2rZLRhQeIkqfK+Z
qDmrcSBTh9Wb4CLlthi7opcIxS7PFO+nWHg/jpGvg4od8hB2FyeK7bxgG20i0Opd
aA5n1CEOl70MXSpe/pXC8h8uSR12YN+HGAiUz13Y8pkrQccPhCa38N51Letm4j7i
M0U6kNWMBgsKdT7vvUdntvW7APJsOT+xxqwjTi2vSVfj+CxOWChdgosYO14dslA3
+L9sy70M7edix23WYKAfigMPJB4ElQ1VFI+EwrqgTLZevY5rCVCXom21AM0lKAH4
wjcGSgTEtPktE6FJs07+xsIDL87DLYVsS2etZzLoFQfLIm6uXe/nM983B2B46HFm
0kt3YvkttVEaE0hIUwh6kiGQf1aiiM9JjIJ9EqJP8a9Ryl9GxUhGD+kNza5j8q6H
rF7hiSSG/lgbqQA7WAzmjGIfvqzs2OPB2Zd3l98WfxNOucC52elwShSJP/cWrEnM
WgkLcj8ZvDJXCeJ8PVw3iZz26LO+ZuNbll7HwZ096xEiIcXw7wBK4EM4UrsMaOFk
NOGW0hSZndRZMpUkPCLbpkq2txb0ZB/E+a1l2PfFz3Hoj4XlvPki4lFSxHiGyF0J
3yNNn57GrUEtG/hh2uiaVeGlxZaeffeUXy3ll7xxRAjEGkocmAbloh353z+MEfWT
SJmZHiMC4BmdHadGpooaEFMvQ+1w0egKaJC7PqDch6wSlgWYOXAMzAs9bL0U9lhJ
6xwUj3SDCWxyky0tZnOHv9D/u6/eH0k8P3CkrhQuse2aFBvunbUVsiy957NKLhGh
LVAF7ANxcs5f8EWmzTyW21NmtRymZu1tdqkO25godCbUHc8dN8CxPgVBOVuQYVhp
C03FK9434YjmOlzwfnd6g/Nr5xRQQFZ7Qaz2jMy39YhCn+lsg4zHTARYg5uVdxDq
eNZsAqXUquTvKusjNoOs0BIU+UqZb4XTButCuYPDBNNH30DoV0fj+a+yB+eo//bq
UoR6I8JRxgVzhmVykb+s0jJrlBriARvppSBuzDXS3iijlflny6FKxi/CIDGFeklX
wZ9i0mNVKz1dDvJIvD0H8QGeEKlyGBL5B9FONg5MOxldMex6IBcI78JhR/aEDM1Y
shzsQksW4S9QYha933DVcRiNYWikRa8K80jj0CHjULPeTqCkMN0/F7sTCj0/V0wo
/Yh9VnBFPidDbsT5qwAhUFd3gaaoHn+c0342kswMUdWftjKy9JuFQBHg3pt+E0jd
qH2UUXhhSn8hVMehWbXU1U/BVSffrUmkG7crn24WPaRGwSOKKjjf8u/hNdUaPg66
04lq6Bq6tDz79Vp7VgbJbER6HKCk4SnCJxNyiMExxCI1WEDaqZjKPJEW8GaGjibH
V72Btoq2FZ3BEVvdKsClrfx7UCVXldzSb2C6DEd+cJt+w4iBCarGBZmCDEJKpZCu
eEtoszW/HWEQQXzH+kyDZsGWzkLFOe+1PIgTuU13xFfoVqK0lJGnu3JTqIetp5G4
E9cUlb83gPqZVnOIU3iUYazcCiyjso/NoZ8uXaDDzD32XPhztuOsLVTO1C4qt16F
xrCoKHypvu59KZQZfmTOGv9mTlNFgr9SBidN9m412e0+48BaEyLZloxCOU6x3uug
S0juzcuZwMvvzTl//lxP1+D4zcSqxVFI7It9YfIPUT52lJ7J3DyZBficuthXp6m6
6XmAQOuRm/ic44oNOv0N0/1JmQAKekdhuJDiWhxr/dxMSu+7v6ibP5L3uLnwpGT6
YbnIQYe8Q7jCMWiKr8tFhENO2x722rvbpCLhmGZlCHUJvvQsSCJx5sfQbMhoiYdQ
naX7l2OnbidX5YCDK2Wpjf2nCbYpQ8bQFxmKcJ/qKOWuxIPJFmKQQHIaT0f7YOmP
9SwomN7k96zwNTXl0DSKQ0FboaeNMiGsXOqDSI4sUE9PEKfofERX1svIf8DuKrDK
gjDgP3LJAZpWE93OU8afupTYoHrbQaDd3n0IU3iogOzKnhrPHQtk5/TDnDr0zzH6
yFOOOeU2aWyC7XGB5kXRI/900hQ/A+EOYrQqUlUGVcv5JUM/b7ROu23+agXFR3WP
Ar4vVsCuxJs6usRz61Jjdun+acuLHuiirE8SAm3Z9xJGbJlZNXlPLoFd7/pMDMrh
SDiV+14fxlyhtSkElVFS7+JWiByxlo7HADK8TO/c2mefQhqOFtHeNN5icYqdpXRM
FbEmv4BklQp60JCn1fXYG/URD8Ex0vdjYVmehifeS7LvPouwvVwwg+6zdL4sWmuO
wIxGW6hloTgwx6Oeue9dvFXnPxhvVy//IknCuZ3s+q/Vw8yGKF1ygITIqay92rjW
8Hv1kSjLJl5QzmtWNy0P253fzbdaaIsiPth7hZlt9RWAr61mfxB/4muGcBlGFN5z
NLAI151zGtbWDUMVPn1YTkjoK8onfgwnFw7feN9a7IegNssbysTeIoAZqHNR6AUB
jMTohHtmekhxrZMjOkD4W4374iDQkiD9FHaLZUZWi9j+VSMyKTuiru373wYeaTcd
t9z7XTQtjgKv/HBN+H8gB0QiAw3Q1zYBRqrt/ArPT4gISeaTcAid7Wve+hc0Ub6Z
+5osIvnGBgZgREhl6XidfEzGwzBD3+KCpAaFgKhB19pH19mFfwGi0v6K0/5g0KxM
A+X6TKrhQOMzgm+kH7NQwtvOimEG1DDM9oad6BEROiU/vLU+LrdT0034ZpOeGnxY
8RyH7I2MHLpvqz9eM/CW6NVB4sb4Lmf3bfMjGeqbdU0fEtGeZICfNUiIhGPnY2Oe
qSUxjCRQWOREeNsODx9UchEmC0dvg/szMLhqg5l8j4zrBLTLHh/Q1k2qL3/L/wsn
/5mxcyNk89EN0lFTh/3CaC6fyxlSzIRWHtHFrmd/9Am14hZzt4alT8S+42qrsdZC
hGlttFpk+2hq/bTla1c2DbhCgc95u8zMlPqNTxAwTKcD8iqPWXXqtLRVOYX3D/aE
w+W3tReNe5+DBUO46PlqlD5lPbHLVPAdEfyhPL1xSX/uBBlhSuMSvZwqBVQj5fGP
idALcijoklcEgd5DBOJLTTL4861NCdpQbFc87mOGlEdqr1/+6MNF10h8LjobFZZ7
MZH2SQ6+26hpcCUMb1z/AjIpr5/Y9/Dgrz6S26QhbAKsR2SR5YTjptNxap0N1vDJ
1Qa8kW43C6UIYtJkJH8p2aT5BjwQHw57P7WHrdBR30WWN2tc1MHnR0DwoB5t6XXs
WI7WlM7MegGjEEI5e2ayLcZqyPl3mXpEZDzHJ5bOfdav3C27Yvzhmxa0Q1Zvr1xj
uG6WRJiAwNh5CDk38rX0PqRbsfSFDYalTWk1+7RHtgEPAHXOSjEuUleOWJE2KiGR
cwh3Yqxddw1ECP+iPauxK7ACj81B5MlYyAJ6gKiz36nUzkMZ9oj7r+1ondYAAplV
pur+n3wAdgGGaPfzhPqT6H/phVUqaxhQWefHEzQe5fvaTizlOez/fHTP2wO/GZJZ
oucsNx5lxSaA85dz0Bqu0FJZYwCfhDK8j2xUEJKlrkbJfmw0mNJi4ZcZvuaat1Kv
UMFaCNBONtuyGWSZRN5O7EuuY5li+ltmvXvg3OIlHdyzJ+1SlcAkrsoarwEzcfnr
YfcqL1OTDW8ky3a0IvyZe4GVRnQxHcQy0JGfrwPMYJx+n7o5X0J2jTlKfiHkSk7r
BzbvjOmAWZFyCtRrFRsZm7xxQtaX0IhJiC53EvocW/PPFUlC5ZCaf+Ih5XW2kiQm
V5wSsDk+uKhLDUO8sd1gZjt2JzSMdYWTfNsuNrhXpbLDNCv8ycF5qEvNfljjIf/7
eHWLsYrQQA5jxwvT7rwJPvLX1Enoj0DlNHSqXSlqgY304vgh6hz6Bqp/yoLMFqPZ
FyOHiECgE0zrsRnf+g9XwDbW18td+tRwnRUGxxoC4DQgoB+3g5sEr546YvZmqv6P
vZYBFRBN0B5SttTi5niBvbylzDWe1399O2RfOqO7Jff00lG+SG0K/enFqQIEsszf
zYJPOXE0dSZVeXpy8MXeH3PerlYPpXuM67gf53zomNzDgXWsIUjUPzZfYdyieeAs
3cQAdLDjDNqIzS6KKPlijs+/0GLkjbtvK/NHUN/s6XI5okOviKvmehHX5e5qHcaA
F8lxzRIhybxwyNaS2DuVyj3aL4WlzPzH9CIZ2kYjofhFRJLQDoqtUPP7ha5Bkcm+
KM7jjrRPO2N8oE2Odouve6lTjJLZDTAC8W6YFeXmlquFyJh/pgBI3cVSRtgxYiwV
LSB28frvz24y4ZJfQOxRc3cxI/ySxzg1C2jC3uz/XBKDp4kBvkuSNHNmAW9ujpEz
3aiu87BZpNTAnLW/ZJi9HdST1DWcemjIJu6YnWgvRWNE8S5hyP3vkGYLnSW0MK34
nrt5w9ghUnefY0TnEbRS6+FV24s2zWzmzgO5o3xjI95jJ7TcuAiwYLA8sIH43Idf
hylzNfUQ3x6StcDQbq61PZfUmKRSKpijP5U7JI3wudwQBQd2+eZcwiMkAiAV4XvS
tqWAeGIei1w4Z1NrOxKI34JQa9ZpMXRG7UyHtJUSS/9e7VPcm2tn3BJ0xibYnl6s
/ILRsiGcRLIAb1e0dENHfmUL6o4WLaFGLFAM3fBAcQ0IF9WaQeHx+d5MMy9S9JyT
37ZTEWSTeJEf2phzwFmtjuK/7QXqbfWP9H5JWArXyC12fujjkErP58e3n3bmoe1r
0g2QQ8XFWXdByDmL1Kv2eDY+eW9qZDAan0l4HnXHUa6jtvauEctZXzdwf2fxeejy
xTDN3DuiON0cblRRWtHapYRTIgRvWR5zEkpQl1NBjd9GWtUklXQcpqVM8FLshNGg
LUWAqKOK3dYlotaksw+/ZzQyMIA5RJQv/i6Kgkq/ZCh3AVK4XF8CzPmsOSxmUUWF
/twglDrQguGHaHxV+GhZPyFBiyaSlAP4+7WUNu0AZUlE/+qwSI8AuOem6wzryPDW
TGwRe0Kqmymk7IAScqCmVQOjjn+jxiaof5TqJMLf+4kU+CDOG22juAlGcZJnTIJq
39BE7eaEx277G+Ci15BehSPoW2axYn+b7jjr5mSnTkrCWkRiffJsOM5PtNWNBiA5
zGIRFTMqooQoxeYm5vzIIdGblC64fgzkiPBnX6bNIU3vzI9h1RoMdKEp+GPxfl8P
rBWS5iPE2ySnmTkMXMARijpSho1sGXV4Lx3NnzwbrZN5dpRc7gIbzTGLsFXbU7SB
sOS0FJcS384YwJPBfDGm3uOTHgLaZFHIwqOyyx5ZXrZCZzIrAAO0PG1tiyhdh3NO
EjlDcHsORRx+hxPOeoWSg5fUDHksLye98qsvVt7ai4CKHehC4C/QhIOJVlOrwueS
f/paGnlJY2rVTjIkaJpMnYKARAPfBJiL8h4/M7rfTvoUSGeKtUgFQ1z7b/l+0PX8
QOLBhpy7djocLPkpssu6keJy+U6pchmrhQkGGkVqUlCSFabragctksFF1yT52exB
4dRVgWV+TyisLxqIC6jAkMJFXLdAx3ATz3dYcBRPNEL0lmx29/U3+Dpiz4tzfRiw
654pDdu4mVMfF91VnYtvekCLOTQxVbrT+fKXGBLKxBo1dHyiycJdciGmNeqNxAL6
7UN3zRJMtxMOlIVMU//OJejYSe8FYQVDs///xhWlhJx/kBaEPzWcdLAOpyybbIgG
ngbccy6+jss4uNSgCGYgYCatmCZAYxQZis3qrhE0RVMAc9j5OLbXPeG+tJmIWnRm
YA+dx5FtMr3wWgK5lzDY50EEEbGXNR+O/MhEOad1jT/25DitFUI4HY7Mw5vv9Sy2
c5ZHIgMCSrYU7FRGkDSYF4aB4y/KLD6I+3gTR0IirUeMstSSX3VaLXTVKExd+TjZ
ICELNOr+PN6bOMIezAsU8QeQglGASfrrWN6fmSRVDNqBcxVnApogSRz6T89qDYrT
OjhiK7H83wIRbQ7+gcMOBmPiIcvSfeUeZFV+olz1w39HlwiRlMFFnSKBu47LT4dA
txosi27YHv0PTJp5di9A37p42gSStWmyjIXjmHUqx7afnmG4zWlP3/UyuA9A4zsV
C0SWaI2GX7XTDHxevMgw8IHG5VTVxzFfZftzhlfyQkrQc+hxwgLXEjVQHbf18vm8
41tHdEtTsN7bBiy4K5wEQ2DdyNJ03cMKFwkJVbxKh4HFOBM8R/hqwn0TINnrESZs
gjnhlIiFNrmso4HIvhU3lcFXMYdXEtz0b36j+3Z/G49D/n1AIdqag2k7DuRCrPed
gHteqC3+LSHV6whpUSGSsIa9o3+ToRvNDQKxUKZ/iEik2iksb8s/sbsKPUsYrlSx
S/de5cxnttnICk1+ayrRgWE7q9MqzFjDwmFgNQ+JtgFheUu+OYqJy32n+bIA74R2
fo9OKSRgzZLn1VaNCQ+QE/nwqio0bdM0g0vMrxCF4C3mun0wg7e+QsabQrYVzKlv
0K4vHzJBTu7aP7UI945VAKn4coM8oef6MRJqT9j6UVaRsPp/3DAY49Zmh8Ai9ldb
epW0hH7LZorxuhX167odhsfFjunq1BHjDGTnIcpxCRL2Fps+/5Vd+tdEiJ8YI+ZA
FVe7ggR6zX7Mhky3LM0gKAr3Rv84Nqnci3IsQeT/EuukvLzmxaFYuWbtCXOAaOyK
jqtjmW/YSgnhyWi5hfz3u42fs2La22W2LG1mqTqtK7SwqaW+KtYDhDZJQqNfDzyB
QD4/opAh8GJWZRHWYFIgcFtscOmy/oqyqyWHC/Zftw42Zjq8KAQIvjnrzpswAXgh
/ULDsjQW37CfchWO4SVm3fOiS+nUXuYeAnlupV4xMSqQ/Ynv3q/XMrXl8NNXLy53
bpUxPop7GEQR5H9bd+AJ74D7MTysowAr+k2Wtr06DyZOUP5s7Y86VX82lC+E6Cz+
WBK7AU4mJfFaqI+KZiwXIP7WkrovRXeSZ/JnvPOfB9ikBYXj5SDS0ryc/wJUfxDq
XITelU+Ar5FoyBCf3bMMggSBXdC1KGF1JI8DyW+PanFhMLiCOJ7eOoqPoPt+692o
C2XYM7DkyHLbO4D42L56d2N+ssDpztH/GUmGsx+3s2Tmwrb5z2BOMJ4IAMJMM1kN
br3/qa041SrJXxXYTqWB7MoxmBfaqOuHGT174JhLWrFz3COrHY8OMZV1252MexTS
N1cl+knHg9i2sqjeu86HGhSRz2k10sOxbFqIOQh2v0y9WV3MVFRMjEnctOuHiVM0
8N4RgCQ2Z+Mkdgplnr5C+sGsdwWv6cLtLphtEYKJ0DX/K+pSbJsJUYdAfhaCF+4g
1RQFmCAgOzonMweVmv2Tol6tmZ2v7kjqzuj9vsykpYZNk0/d1YCf2hu0WKC5++c/
VtkV9HMebXrH6evubhtQtF3yw1hR2a/Mamidx4R6FIYk11vn+h6gR2sltQoilF1s
9BIUQxq7CUsXTOttIlNSf7Sm29HejT8lbky89KtZ5jn3yO52OoLv3Kq3NyA5rxVK
OTnU+LbM6Zk4G9dMQAsCHokmB9AiE5dELOTHdGPUyw9yGNHTL4siHFPsHUiCDh4N
Xpm+zA1m7Y8F3Su2Vqh5TP0NNTkD7RIfWEcx+djhvZU2fr/p7oGZhUzUtTdFJPd3
eCp5HrEQM5yF67bOe3VPnWcLG5CjVLQ0KtOa1RzbFS0iaO2y9NDc8Ku47w6iidxx
LPMtCyBMe5tWeDy7tc/ynMbL9J4YPGgSJTd8fki53tRjDDOraIkN/a5KgXc4PFjy
/uEKXgpjM/dfd4vWToBdd0gLYNk8Oyc5PjEPQj8GNlyt67VFbV0ds6qpDGak5SIh
2ODe1bbquuv/Bh3nzYlxMtdbVexrSvNdAqzzMI3dLGyv4DTh75g5aQiEtspNYMeQ
GlHWF0W7yKIFu3xnrAzYoi1On3heubidf0s9jetmrUat+gdk0i3qYl7CYtMdW5UK
FF8k4ZMjgJg63kogLKWmJPefY7mbFIqHbAPw/pWTQKOayCazxfzutU/EOqt/dGlQ
Aadw8u3ilWzGn36kVMYvnYJfnDMUUEnFneeyMgnFQwnsA2TvcJJhgSOJF53SQdau
spwIwnAbiFpt9nGATZt4+zX7Cx+kxv7LJnKbixN3+pl7c37i8di/eu6kDkYWzuCm
6dOWhL8DiexYsJAVt0qhgrHjaduhfbkH9xUGNQWK0YD4Om57WVZcn3AbB/yUYSSr
FXsi0nyM+WhEr4Fo/v9WXz8GMqs3hAj5vjAxBaAMUJCi6nPlcXH2Sw83cppVRBkR
wkcYFX6y4KvggaUmg0o+PqTH8OFlLHD6KF91IKYQSpwa47Azk7MtZl0D/VDWMOvL
+P+4F9QaMD9lLLBTuImSvPsaUzTxVIffIUoFgi/1VfMFPSrpRUUs2/+R89LrSIIE
beqw2om+IZMN5vn2aKZqGOeT/9IX2R2ccDspkF/cbFqH+l3MKwuIKVOolUAFRjsY
HVuASCz+GH1H0lNJhxgJXUkYg1wS57OkNl2/0AvyYNOabDCODABJ3D6BR5gjyml6
IB9HyGd1FPCWYtq+/H/TvJEgQXGqzuQdX0WcJ9GsjWIki3CsG1+np/6M+Z2libRV
wtP15gSXkg7D92hIPwT0bCjTcRzYfFLezcZYw/5p9L9X802NuX2OekEuxKCR8OeB
42t7VB+uSFI3K5qrqrob6YFjuAAYK8wMFAiyfeuS7ti2b9gvLyvt8+wD5nbakx84
aywAipeO3MvoaKL8pyDzX0CQH5GTXtXjmulEJ1HTZbasoAFr9j/rCA89LAV/0Jer
zREuQlYJAJpX4CthaocY2BomfDuyqwadeB421NN/qtNianZYsaeAx/d56scmjTyG
CRYM/yvvKkTPVGqPjupzzCldVjfwGd/r40MBQwHMQbdk4e/QG3eqYw76T0iwmSS1
YGXgu+I1xAU8skfARIv+2IiZDI6es1H2rpaIp2Sp6KDxXD5MaL2Ukf/+/MKBTL0f
Uk03IX7+aWzq58zuHZzffpFRcXqU5QouEdylfaPxfegdL8yOmRqrfuGhWw/znMpx
11LvrXHkhcFzqN1s5f0JDGehH11PFMKWP+bNcQTzpQbsnMhsU0LvrvRkZO0L9HVh
4swzMgzM98Su66AekkFwed2ULnSpdD2IG+l+r9hsK1EWliEMMUt+F8Lols8G1Xgg
04QgA3t0xZ7H8z81B1ooIS+WVu3F54iBvAzQZl3TXvvc8LNBfpunYUtRhDnPwowI
yJR8QvLiVoZSY5tbnDa9MMkSvjmACTroEmFDw2qVKsqvtyX4LgA914SfByOb7YFc
NefwrheGexwi7g/m8EuIZB1h5r2dtB+skoyUt0weQFjp/1Grqd3U8arOt8WaaF5t
iX2x3Yi/j6sfqJyY5l+65Cgz55kh/OGSOB6dGetcypoEH6Jyntqn9GULkd60+t8L
+QBGws4mlf073GRXkC0KXUrCMpU8kFCPUDoLZBiaSQab9qH4GRIhxPSf+LVgHyN1
LvL+AnAE+PATHbrzZhdd1lA1yvSepA2MnwYJHPS8Q/iARcxzC70Ay/AcFvxqYXns
Vpv4/fRP41mH93+j3yTbdjkN00JFNatkZsv8ParS9KjpbDP45CtUypy6EKos2JwB
+akA/zMdaySOnRBOHMdUBXusfEm8aTDIoYHvR2cMV1+dkPdz+L8NUcy9knJ/mTnk
JPm+afmF9m+ES1UXcv9DFtDaFkrWaKvhGaVIxJx2awBlUcS6a8K/n4BiwBeJlv17
Qz+o3H49hRSdpfHVRL+E4dVbtcGD5I7DhnqivOi43T01/ihKmf+Cz84bwr7ARF43
lQBlbKmhHFpCtNhgjpaulhGHCy5yfiShgc52AJyF32gXRsPe7rwD+0o+EhMr34EE
+QfuoGDKMCv7uRRNs8zqGOVQQIpP3x6EaU4fPDRld9y/AE2nYdSE2uNw0mvqBDI7
0kS5E9QhkcWSB4Qf3p+9SeWDDuoVMxrYtOOiBaU+SI5lVJTAEpIV3twTfvNPpZ4T
RaHbUKkBnPqk2yqFMrdups801YFStErNLQj7v3uOKrkOZJGDnPYoW8zuQFVM0VjC
krwm1ZYdaPfITO+4DYl4kgEPXcQVTSQEhQclXFWnSbGzE0Q7AQQePshvmVr7B+/d
dUf9LMPZlHyV/7EwrpUkwjae/LZgcvoPBiRMhlnkorvz+H+HCxgCyDskeOX+XVIG
Zl55V3d25qUmflE87gJXdJ1ejk+xG9lKZFch7CP/EKchrKcehyw98M7jGgAA6qFX
W+Aw7m2fuDalDPGzkE6U39ixNNioqWQglUJLoST2DbK6UfKpEUbNaC3lDXB61uok
G+fXAQqrn+6Xw7N0e6cKPxmQnH275nKiBMjCht3fbS+Q0m3SwE4zzzQ+8synZMkk
FJbtJcaeiKCgMV983gv7eJHPenB9aCAs24sHRlg4gevH0jAyfZfD5O0Sdn+hCIUO
JdqOPMVAMsXm6maR/PjOFH+tSCem+Nb9Rgg08/XLY+pN6pvVtxFIJO+hkly1QdJW
9WM1tpsa2YO+IKRxiuPiflIsXKqb1ooNPbgnZDtgqtmFtnlzHUaNPC6rhQuPgaD8
Ei8ubmVhLRC7J3b/OnHlA85gipkv9lbuajphijDhGl2tZTZDJNIoKha1x1TN3EHl
ZDlMiCsg+S/Q9Q84RfYI07OepcHYHYRX9T8UWBXDOHnQ/aYe6KHI2SCqlKsNXeAw
zgZkCqvozTv52rDZpS12dWVGWTKPmEytNOkOWOu1DXORpL/JWwVdIwkZ878VwPbT
5CEcwJsXBZ0HWIJF99A9T/modWQ7wczHGzYtqoPfnKAbFBDYb9JKrqiH0Mt1CrXa
B3A4FWPIdqD/4t4knxGac65+16Y9yVHUAeqjljtN+hMY04gC4QoN1Y9FiZ2UIl6l
len9jT00kBmMQ6H8T4Xg7+9+gy2Cm4zVLWjLyPQB31kLfsT1nkrGFOH5vlbFcelL
k8mTCTkgMHiH9Q110Hyj2CY12urzj4yVlh5G+aKfqK//eFsiTjQbYQRzJffFKFaB
AzjB1as/WqXQQsfGEO7bHxj3gVNenRDi46ob6iRLGuYE+l/CpIg/F5T2u4YxXcSv
v93VSGw0Nu/2vHJ+CBpL4ST+azTYddDmo6Kvi9TqI2WYvu0rinDkIaUgnbmd71ml
bWa0voUmZHx7opyKtgZKSRaZBfShR1kb3++xTo4u10dlZGJnPIbDfxL2nAd5ZU9w
51SX3kvGvqb06TxQjPNucSQcBYT+Y7he5694ONtl4S51P5a2sE+MLSeezxuycFyZ
Dc++v70YARMbIvwW8Z0unXYwHrKBStPPSPi5vokL7mim5jQzLpUQw2v9i+KeRBRr
XWTcnPjWVu9pC16EDO44PKp7LFhJyiVZ1Rq/MeX31cR/waPGxFzLYGAb0+vSIh7b
2aNUPX/5rfObRaOMGsB5Xo1p1YqVBMq4OZuWTzH+eHsrXGb7KG6AcK7y/wXhgTCW
o/8Kee2Z4I0vE1ziMd2WBbtqoFOlISEzSEerAizuE1u4JUhKTkF4w5jYHSBRqBNO
3ARKEnvhhK2TbkmH9QuCZ9mxtDmfCySv9yMbbcoaVEFEtrm/Mha6pesX8dIA4Ms0
73eQLEPPS8ax/c/LYgx78y4Oe0LN8GbA1LhVN5R6Kv34gMU71qpaCA4OdccITw/8
YoIBOQcieXzBzvG3hpDcW/E2XHzd4dN1mCdHWaVA9/6j7c0t9kAmKqsVRDlEgZ4n
p3453diVRztimoNE6ek2R38PbaFyaomZkH4D+wl8tLJ/Nh4WTvZpCrM3fZ9F/N95
nuLZW0m+HkEoMjFmW2Ks1ngG3oWoEWWWZ0jN991adgtjBWFg91BxfLxsBuWnGfqM
sLM/UDjAAA+aU/wCDEfj3dThPkuLYBuRqFVuT+G84jlOVtjmd5yw86C/QxqAPVFu
NfePP3hStsFPyIEcsSRu3qoobdHdFcX4WIdSjJ9O4Ag8DOAKmYsWz4unDNy4Fthi
jxRB0iEv/R2So9eJOsZVqnmDLwybE2dyFDMVHxmBzki04W6KqlFG7AB6X/DNroy3
0bisO+ClD8n2enWf0p8Aw3/M8xxbZxrVRIfmgtyJ7GFXjpQPMSWg40l1UZpIj/2t
L3a63tHllouwd1/vAjmBL7LSS/UzFqgRtMJ+0mJKFCakplOQV8NDPxnaGetSsw2v
+84ov9WnchndAUFvrg6cNSd+vAEKQlTMTM0rUkjRbn4c5QCTHyKDiRBrOnIk4sKE
UTj49aeQ7CUPzpxHSpOP+9ug0ZyoVa2CeyuWdPdV6O3SrplBipNVchdL4eVM4qve
5B3EhxpKc8KE4msccfuaaDjOQP+JZ0FodXpgPb11g0+zaIb3eLv5BRzhJGGPApuH
anQ7nwmkI2YivgD+UeDGKA3IX3dmnkCmmPuiQwM7dxA+DHlD+88QDI1ic1LL+AbZ
AGOKLjEAQaAaI9LblOAwiE/TqrpReJGzMpt62v9Z9hxqX9+TGSeg/cCn29d+8o7f
mDz6WeyhO28G5cxB3Bgn36CTAG3C7T2oaf3wEqbIcBMwoVeL5yFHu8Z/QOJJScFk
clK1A3UfYWU72RPzZTKfnYTkOOtgeCpkMVrSsE55MYlcGViVJbVXNUR8XdmP7iY8
vY9tQ20EH+tpB2vB3ZwXlzeGFbiHiRcgX8T/Q/WvTsC6h13Q4B1oJhjEqr5Rwbp0
etlwffcs5o8R7OnGzOrAn481nJVSbkfJ8AeDeakM306QIhwfY4a1d8ErmnQDSsg0
HAQuZbMA+k0Mm3oMyKeBxd1vVx7dJPC9o5BjFl3BtThPJVlSHc0cnJ4gpuY+6Cx1
qqvEK61XFcpRGRMsC1+hXnAAJ1Z/+muZyuCDBWYwg1UkxvllGKEvYFyCESFpwEWk
ULb9WuEb8KnA0iXRlEENHg5xszJsn3MnaKt/qJ4woQSSfDLSpAbfR7JoAJmXXjtP
ORqSCSIe30o9gV9uEwq9pNdyzX/akfjpwiY1hUtiY4H2/rZ2nc3JNCJILH/uey/r
+84vkxKcSNNRFH9kfJvIARMluIMRfe409k44CY9MGMrTVsw2evlbqRkC1UY/XN5h
XOYMfOgccERWR+slyU/nAnO0132DegeLD3tKXB3fwM3rGSkrUdEIU3vH8FuXKEqI
4txFppwbH58rIexMrNbCtjN7requ2JiqAuRDgTfEDCVRp5UJO92NrZSBKjg+s3TA
llowjlrG0BOFLOnyVc5zW6648ZgqkQnduTPAML5v6/9K9GPeGDr9WZ/XGFr9u9nk
ItbDeVo4W9/JWSHEOpwQBmhA6zNCMcs9ENPGvf4GsGqvfBPjzkm+f9tPAwNZqxt+
hpXSu+9L0gxJIKupdrWUkSJj23IIy0j36+ei3bwKMHKZUYL7bmcPZuhAvyabtS2b
aU0fT2R49j/0++VJrgLcLbmm7ZUL8MYGYJuL7Znl6hNWuvIzNba8mBu9KAWCJgTt
3N3Cjjq7kCDEIvS3rQju7mgrK0+JciG3h1NKqi4zV+NYhoBUACb41EaZ/rl5vnQU
WLhmXwQHnUFLpuNWMC7Iyq58E/PrK1PA7L5uCJmoalNH8CEUn6jEEsUjYK0qLV+O
V29vWQLNJotFy51S024gRle1oUwufh+yqC4q4LYwTbDCUOeMNAit7lCWixullfOH
C1eyKU4RrgFnXgySfltVgjz1c9Yo3cG8H9fTSxLoHiDm0Ae1OwyifHZBTL02y55y
vx0+/CiLYPrjjdxwb9p1LZ6zVyxXew35r7G4C3ePZE0PPj4+3P07JxyTvokNIMwi
BmP+PTAg4jtUFawWRqS/ozqsDw0Fw82+ZHnQi0oUpLOOnyIYkW8n0LkoPAc8C5tJ
IW75CDZQRtEwfILcbAu/xY7JQ9f7cQlRv73CZuVcA8y97fdXmefFs5nVUpNlY0R0
stqFLV23ZsTM7l6XnJGjE3TWSYXUSWmV/1ZhEN7zMoIpWsFHewMBGVi2wRrV8Lmj
0F+ZkyjE9GApJi4WEiM/vevS52ep4CaTFj8MEcKxvwlfJlQOFQXOXXaoPEBQwAnB
UhcZuZ0I/2aKszkA5Hcqj+oOk4TI90HrwgbZiZe36OG3IjpMbis8Wx0v6Q7knYZ9
8O9F+nLJA9OfFo7wTLL3a1wTA1p09ffEPtu5e9IElZbXNTJHS+tLk3XUau+HUF7O
4DAnDYCSTJlFhaxfDtHaosjCihHc43LdbRIU5+LPIGELGvkz5UZD4wniPR1epoLJ
6n/QKc5Vp4vTLpfLlCQH6m2Si/ehvIO5DTDu9fYy85bKbJpb/cMBaXhgjZDmXsdc
5/QCEyE+xFjYtzDIPSaG6NKmdyHGtOohilmLkstWm75LEUUrbAJrjaJgiE/tabo+
w5RuCa329iVkP9cK7Tnv61wynUpnC8kO33Mi8hsB40YN5nntaJ+77kVJH90cm8K5
95zIwngPA2s78yrdem9RFnYW8dItaDiKtfEvZv6fhyvvPG/MDvpHK4GMD5oC8XSs
37beXqhBHI/6S6au8UAUL7PFqeuwLcFrPfyjIq2Yg5ecMaFnP5KNqI58ZV23qPRp
3Zfbjy56FR5mzZ8oaXraomixBIn4yu5kjMTMl9CBWP8kMdr2CyKfcgjA+2J+PBZG
27vUog08oig61eY5KgnoMdxTSPKj53h4aA1r/F0ikRnZURv2Ds6taBnvsBLwfnvm
K7/D2rLJFRqaoAts+wAvOZkjZqm5lJ3phSbtGevp51oXtANftp9FuGHokc8JxUJ0
e/HJZRBXLIXfQbkaV3Xe04TbQIaeWoxP1zkEXWksgRN4Ytvxn20Ju7xD7DmGSwWm
TjYulf3vU6qgFyzZHSLsjm0rQIgRw/WWbTGzSu+FTqro3f657RxcTXjlLppIc+p2
H3uJrDdYsvH7O1Km6vHIpT8af6wNokF1Ayt5LO1nxDWwIBp7pSd/JsjuLhT3oLc2
lIBjX8rMT4WGqc2BF3gcK9/0TSz1MOGy0TyBO2ub4TnGHu6/r/Mu34xTBfV7T0K6
9hwltCoiSJIrQ2Fn7SG3qOsf8LQEK6i3HDHymRf8Cxs7FIs+7z87OS4lGin/cyYW
7O13fr7velF4Ny/1E5wcZkQEnw41xjvYJRP4MFAE9xjZ4q0/TB9sR5huijxfj3gY
/yQM6u7SZheyar2DF74tYJkxOgygHqjRCDgIAa5IaUotS2pKCbk8q+X/5hNTsrxo
JssmHVMN2p5vQfH4byRXTyb/oXM+b2deZo1w7rHK8FGjS6mNMuzL5uLvnw+ADmu0
gsBNegzVNnxU6nKZmN8AoSF6uzcI6xeNNnZK+6tmILjrs5RKCS/5UDF55Z5olw6e
mMQJvl0fpMh1q2lx/Hg/Y2GXN1y1T7Ihg/1CIprVes/EXUcNKhbF1GxmsQxuaRH2
bqQ6LAzq9X0PhKa5M+KPeAWk+w3qAXCUYH5u6xvc74XDWlKGxnWUKmAGSnRUVUD6
tqgNDsm4S9UllZVeL6QbxX+PH5PDCFljqEC/ZSN5TMZstj5DUTJxt2eg2agP8AyS
Xjd6r7pn1xq/jMORq9rf9ncGtIp1/M+q8ezqpEAyJ4CRzkzFqtfRalvM4E+1VGRK
Yh9qYUctjZTzTp0OF67UGk6rdh5FZdUNujpQuhb1gOdZKsBsPkMZ9343j8/wUsJB
MmLmUUitS4pgnz70Szj9H+cuKI6pFT6QVWLIBT7CmYAPbT0WUFAuGvSGbjTwcN75
Ye2TqZCVScns3AJWErEEZYZYQkyX6EZ2CKaKEWGo7tOPYPXALzOtHeMFpT8xBO0m
bQkD8wHxSTd8I7WlN1/6+C6We7nqaJRufDzX7Z+Ang1cB2wgHr9apScBxtBYiuYo
+j85dZRncRY2+v4ZPpvVdWufYDzV0Kmmps/LsownPoxMwbtWh2BIaFUr8zp3wHJY
xN9+gyv2sS8i7QTX/c8ZcKjsi4chZO+ow3bUYbvTeVoXOcfHVjosA3iuHB1d5kV9
bQ1bD5HTP/EawAJsR//F5n/ZiunmChwEr5Nk1cLRFSWxF3A7TdBnEoBUd4gAnbt2
Hk1BfsP4ERHOEHvGpCKzz5Plqv+nYHhme9ZLKJZbjZkNgdZ1Ny0LUf3aNPWJNdpc
DxWd1ghAl5Hu6I2yRAJAY3HOSIyTMNZYhoZ11a7+Nf2f7dSwJgPwtzQKj+DaBP6V
93rtXiecvaunofsX3DcBRfG5wUeZHPIC+rr2mMFrznGL4CrE5EwoZaC0nEnGuxsp
wlt2AqLntQ+p9zSLD/PvAWX/hRyGtBvjQQOITzmkMtupTU15hPSPIieVI8X+i/lT
p4rqwZjoj7I5Zt+u27A+tBbyi9TBtnlI97i71vPpZeneX86qwBZOvoLSm+K+5G3N
CyxXOCIaxi8QiL1kyn2rAzP+Ztny7ync/hJWIlIE5IvyD0ejBkg8kkQJUgvoy2f4
nkU86E1MgW436qaOw7todDbEoM6pNIrScpNudGqye3wWN/e/vS4dj87Pb6xFraTz
bBX0RRU+a07ZUs8vPP23l8lsWFN4xdZB0YppCypvhShHWvtVfUGlTWGUU/IkHdLu
yUvJxw+G0JLrXmLAlGWH/O7I+WrAYtgwUiQZnkXrARFnbnNeIea0VjenDFM0NdSm
SH3ETWgNKCsKq4+rogc2BbTEculo/55oDArHQh4k9Z+heuIlTPuCxdfYgJ4JNwyv
yRmEkg+LXlq30NHGVcsJ/QN/Br+olgdl1a7iFYupKAnp/5d7o0MMSWl8wkz1Ejd8
KXs56ALAzX2aFR/7GBTLFlRbrLkIZERNbr8QlG/Mf7Iev5bv6bHmnt3B1i3nTTKs
j+J4JdfdB2xa9Z4ofpV3JPG4Dw/ECvLm7Ei/Xh0yfGOAoPykSOqYSfFdp0cjGeVq
6HP7Pl9heuflqugpD606Giv6nhPQuLwOBlfVZ1/aMtp0OOaQA2orhr4iFUq6uWvt
06Bon1pC8/wSDX8ff1ckNM4AFZC0mBBqis0/S+7swL94fjZYomksSK9z+vPWvCdA
WvSnrqYzU/nKk1EeoFmxLlToLUrwG2FS6Rttiko42jH4Jq5ouEsbnOGr2r98NgtA
5QOCh08Ln3QR2Mz3RAKWb5OpsuDPj5sFWRzbZ8AsLYF4VeVrEY2ftg9vbdJuMLpT
YHRa+gAvlxW1l3OHooXforRRotsdn3VMbkNhPc1mqSKKkh8F2xw5uaCNZRzijKa7
xmw6tYJ12U8K0Z3oFkunNFa7f9TCyMxSZnQGTMUnFQdKFu2C0ExEjhcf7ZNTXndF
fD/T/RbmNweezoFg4pso6fY1rZoNEbcxvKvL2a2rqaj19qmZnIOGoGvJLJzB8giW
Aik7NN9pW9dFi3m9onuL+AQcOhLznNsFhHVedAfdS1FnVxn8Ill1jzA1/dXnSGKh
4Fn454fWeSPWKaqb9gKtxxgJoeMueCsZ/E3qnvRXJghUnpz5dJ8seyg6loaAhvKO
E4Ai0gw/5YaNfHvqOVNWkW9Z1ekcFIVm8BXF+uEl43/EM+GjQbL78LJKNHizOJ5t
I03rXUDypPlMb63sVBfR4tF+oWQ5ChazZ7ghTApuWwr72hqpZN7HN1P2/8FC9uyp
f1vMuyrMEdHqhZvKKSZt1lzK3K41h4kkmJizoPZ2ZcrV30fJhOH5ivI5NIfsr+JT
cc/HodrCY5Hmf7OqM+ASOUBkKCd1T7oSrJ/2NKbWQfe5twGMf7wTcFP7zE7v1xXC
IIzXam6SdIZW5C6ULCj5dW1B1eoHPR1rhKlU2NaAGNqOwJ4Y0+iy/HaVBhmKcF/n
REfo4i5C44FrODZOxWufB6JkwmRxmD8fVZ8CchG0YewMGfD9IJEe2Ez7rox/2sug
01zMqecxBHES/qL+c0tvtsh24O3GbhS94k+a1AMAeBr7If9BRbEB+CaSDdUb5RFF
uOflF3jyF6gAeaFrE5sauFv+g5VJ+A2sM++xARGRjCeZ/tUcpbgl4p2Nto07tXnu
CJlaj7ZjPBJ/xe+HtLtgOFXqCd4/kt9eVOIMWBDJQ21kEWuAVXQkkePz7zQ857UC
URB2zMqosaIhEAf7ZmoVTq5IzCOHuLc2fQZ3/3Ql9O5FIF2BeFDynU/M3v9Jj8V+
68HXgIELDoUFMpvce27C0Am6Nnd+3tS/59N2vMvO34CFZ+evVcxrqGzy97eTjLYp
urnsRX3zSIBAHl7saPaBZfUBA9gMFD5jAIP5vdaU8wY3iAZkNG6dxRwNY2YfHO3G
zz7F0QUQM511EzhDXbsvXlvItaDq/8P0ekwjewlIsVR96Tk/zTpaAp++pvOm02nn
LvN1zwm/z6JqgLtyN4jmQdLiYevh/LvB/LcQeo2CncWY6UXu1r9KH5N43F/f5c22
jEi21F/mpB7F3B/PXbwUcNioSVdmGFWD19G8sUWCZ2yaK/OiV0lT9v7umrrbjMYb
3y+fAyIdlCCYi0QetZ3aGgEv2x4yBWX+BbsyC/4CTLZjZLw3pCUYS2Of7nqLJP6Q
Q5rUd4sfvOIArqyLP1vshPT8S8bojSXZVlAz+doXc443o7cv+B9CesbKE5c7B7Br
GellYwcW/H4B842EBHvYaRqnXknGFIOgDRmqkI40r5XiCGIton5+8Mx3oagFqppB
5+43Mb6XVPNgbs5ZCHMldpsauoQ3JSu1uox2/newnWxMh7BuD1oQe2sNyZYMVtqa
tP14LDpjtH1anhflTsqLn4XUD8X/ZW5E9P3NSyIXOfgG68xiGbkglWbYn594pFqM
5qO23jsZqNS5odwlGaF3EdqZK5eGckovka9DMSuhn9TZieM2Tr7bmbPOdW1KN/HV
wS3Yf+U0SQz19CTBiDdQSveyikmCERJeohjM9F3pouBPIwIC29LRjGvjAhz+UG7J
TuGuRBiUbVJxR3XOx6aeTF2OdD66W4PkZsfa+js6cB25wnTiKkCBH7rmTJudkydQ
2GzaxwYBXTVpY5+A5sCG7dLZWkUYTR3l9xM/XFZkwXm9CX8q02Y9Ohlplkg2xhA/
h27cCsCgxmoYy5O3Kv2Ci1QpTp48FdjA8u8nw+gSAwgIFjkkmPnjPvz8reerOQN8
3zb2txfWGfuej/sDr3oJB28o4GC95GkACHDS+mh8Ec6Ipl3cJ1YC9seOIPWJOL83
xV/l003vBTybxQ4KlP6FbE6vCDqF7AllbGFEqcxKd6ChhRzeb2NhtrMx+6+praIt
Tz7tTDxOC2eCoXrcoHw9JfI+KFKR3a8B9VGJi40C5CbQdodt6fr/+KSS1YdGPzgt
R3hX7O08lWdERpHiR8uVq+3OIP24bRx4mk02UiP01XwlaI7+bOtOFHknXwicuPg8
xmsAeohCOHSLGJ8ykckSsn44KfezeXRst0q0VI4i3J6Mmmlb4042cJgBZMI9YA+a
gzn919mAr/I236V+uF+TAvS8NnoTcKm+FjNEYIHZIYqVzldVF1BllGa1nj2TRToX
j2mVZUKbfmvzMzdenN/iWChOFgcvvUDWRYXjVZFQw5OWzIBRn+BucxKONwc+nZkD
v4IKoQGI2btPyR4zaSLAMrHwnlQfDPKWU1ZitYotX99H16lXyl5VcqQ6WMgPSeVN
LyetLXDdeHVd9hfIIOU8hfyt6lR1scujhvcH6fdrWe7wTcV8ESeN9EGyv7iDG4UN
rHMIySSY0+bT2y4Ul6VLg06Jdc8FidxYJerSvpk0x88jBOmNGgB2HhxNUemTLPKd
bKB7824v5RXMFtOxV1IQRO4+YHcc5kXBZQ34kdM7WujJRq7jBAr0OYmrBmh3atTz
06D1UqokbswZtr4u+KiRhX/z2xoPEByn35T5aXEQs86QtooWqz6qThUOsKPMkjSj
NlK5pFg3PrMklkSingzdYBWZcLWVmlb0JIwNV3lbnWAKGqdQxAwijTij3H3xm81W
jzpr5AuIsHy+BBbB1Qvec6BxR6hOwoBlcq2cbtNySMbXKkLuXvtAqnU+PQCXW1U4
zw8MSVoSJztbdSQbEdSkTWSu6+9PiOON7U385lcXAqqbHHLMdrI1/eTXWuoN3kWE
PowqGn5ephD1WbK0qArGwuLRCbCYln/OIcLuPNr8H9TBZ1lSfYoXYMJ+UiZDP0A0
hpK57BRZIvbc1nGqD+fnoUbWDlvS8okJc8E9e/13GMzkBz4AfWxBjDZjMRSS4loW
DVzkL9AZA5csKchUxodxyMBvLONV3cQwEom2MugGXcZJGpSbVo3UH2w7fWOWwN15
RHRChnxWQSy+TZG7R/Wn6sc3YzYB/OCtqHazNBl+cODDgWcrdQY94rDq3Jwss6c1
WwTAxPXoEU0txHF2ol1LmUUBOSxR3Zkpvcuh7cT8WC1XmNUGJFbO4/oqH8BceTJ6
r9DhKs2gISXJnA5cpmbRycS95Ny9Vx/paKWEWJA5M0jXOX7zc1Gras+AL7pn41V4
ZNJrg60KpzXGM9SKf3Mcrj2Vg5xdwMKVGaShubeNkqPaylbV8emfGRm+eayY3fRZ
GEguZt2Dx6Kwpxbf2f0V7GWPye+0wBhWRjDDWlTJ/t5RD/fp2quLkO0nbVnfcsX1
QAOpigQTi4lJQ/Juh27msVLwhlHkPbfM0qiZAdb9913+VcGtxFKJsjFm6J0h0zaz
j+6cMueaydF+AYBQpVRh47/n36zNqSaLaVFlGKTPxV8Uu76SqUbz+I7GaE8/LrrA
CfOiM6lQC5WTROf/f11DHJ84gJfcsh27Ecegu6ndb9htPhykut9nyQQkoa4LrFue
sVvUHOZKowE0ajf8dTxEYHFQNdQH56KxE04mboafMYuxUFORhuwQjJq+I0ez/REH
ySZGKaxpDKP+5qZtT6+0FlIX1v/GA3nhnQen3M0OhWQVv7gOo1LUTsDvMI3D46EY
y8vDZKqolwrI7K44L3hPqjR6qYwJslXhYb/cD8ONkNC3O6RZi0ZBFcyCBX8YILcw
bkzGTo6MazFKvlkxZygmT7OShuHrmOOpI4NWenKyBU8aUUff2CR3TYSeS3CXFLO1
6sKwiX8ZmOVHDhX1/gWkr4jPkgDg5YU1AeFPIY09zatk2bMJLj5z+8GL/Qjh2CJs
rDTMSyd5ohkRMeKfdBSiQG3k1Bqdr7E5fYyxT3uKAVAc/DOPvz1cvg1AgwUIKpQZ
+PonFb0mSE+lLH0BUVr+OXHVVghtpo4fuQmuKg1Gl2LwnRmQyZ9U2wrQFCaQRFjx
YjB9RHA5Wjfd2D6ycygaS58P1w976s0p2DI8LrUBO7iYeOI23xy57sK2OeL7M9uK
U8NEBWWgW3MVMMEDlMnZI5l8s5gS2kGJQPi+n87wn4dj307YY7UX37KmSPoAg7PD
GtfRkWjCUeq9sRP4if4bB9EqXoqIcJDb4wFXp9KDMkpZ8zYxhGu1zTphHoHUD4PG
k/5NLeLoINeyUnxSiZ+kM/e3R8O3Tp1pdsyiwF703dKR3xyx140caMVlJ2oa2CS9
IjAuUJuuVdbGMqLipaUQOb3testFZC1Q2uvo+vgq/kggSF1jhKdam/vMuw2qYRxb
BESZLpNnbLAZVNfF4J2oCGU6rpZI9Q0QKV+JiZFqsXa7SQD1n1l1x6yt01w87lDf
VAubjCmB96QoAiPY5duRhQOxEEVuCxDnj8hKECu+C0Cby0xoKBW7BHjsnPnoChfV
qil0pjeJrjPi9enAHw99QSsop748ReBjQ2atjiaXtc1+vUwGLgyJB7ezucZ6JPBo
VMtVvcEKxIz7Ze8S72MxnswVjUvGVTWgUPt0OBlYYgrr9zE5RZbcWVKjxqt93eIt
saRbENUUo01NVSc+61xxroUJ1EP4jdKOFp+VOTcDalWapsQFtS8M5KfhhB3zZ7n4
rGz6oAFtiEr8KeQkpsN1S1nG6zPMEvxefxff2HMu6YIZlrkIWGRvXdaj+7wCZkAM
OdF79YRzyZAoS5kqIr2mIfrJZQsUxJiJeFH9v0okAKuMHw2v1UMGRY1+pEFcHbgY
qjf3WrthTbKAJhIewu/6LlKSQ0vBrnfvEk2kt1PD4JqvkZWXOZ9wCS3y7Ve0YhLf
8j5TWrED/MWuovK216iZ+sM0dq1hAhiMVpFck2othZVb69qJDAksLcrAdJUPqhjx
BYc2hRsyo52p/eKR8Uov8PUmjU1iRdyaXB3GAhQ85/PPGoPQYAJEBud6kY+2n5bY
1w/gvS/o/NYUtk2JCpyUGVLnx7j/8uFWUCuQ/ADrtdrLo4t3qeJSWolFWeniav5T
jo7Q1SiLZ2wUEHpaDh3AHBLCzx+jMfGoQXKerhd7UUnzVbNkMkNEtSxih6mC1/wr
YhRfqzeO0OSYWPkB4M0/xIJO/RarxHr3fsq3dfagTq1mwkdycM+3b0/LIkH/YJZc
iQabJTHbKaUkQ31V9NOrc6IqWyQ6EylaKkSlakPscMkMiPSPERVSlY6PbLmevJ6z
QSlxQ7Giq0UMaZPnABJlBlCxN9G/aOT4AwG3L5+toACYdOyHqduBM0bsbq853ZpN
SWWOT7eVbctYtcn9MhGYfinQXFkVgwyyAux9lbSiDOvKYyRGEaOPehLhB/xSn0PD
0CPlXuHZMlKGzGPteiGPBboObmDZOf/prLjbDCRXZDzfoacYPTV7EhqBzxe+fSfl
LkddtlzMrVR3PnCu2NLGR1ebjkmwWt/8b7liRrEwklguHEvPGD3RjH6dhUj+bPvm
M1CJ8+2S5rPrD+Ba+GdYxw9tOPd4Qam6XXFvFWTueT9jyQhVS0dS5DUt2vRZg5Ax
u/XMUnG54UhreKSGCm8H7MvlV1VbZNQpyWg4QOLkXlVH42Wtdrfe6RA4vyD8SrWK
3X21EORMQeFDTGtFeNNRvE+C6+K2vI9nhUxEzS7KbNep6Ckq7EAPyyDIOcnYcIHz
bSY4YgUDsx1of9TqAc/wdjZ+ngnJ6wSvU8dE6oMpATnvVLjNLwVkNPEF/hBwofBX
tdz1RQlgjfD/wAQqwLfIK32Zxq1k8IxSURuER6/6Vp5sqf5W/6E4A46DY9tNSEGd
014kvJ1D2tq7eX3tSTnWFTNfrf0PckBuP8EIVg1Jln8grf0fhuaymErAqv3rNmVJ
uI6pNyVaq2UdLXYtqC4DDXKw+ppaObXiPQOUxTO39OpmbscB818oxgZll8kjMday
8PS6tDhNcIk5yktNryvhV/ItKIaTlH3Pb5/QCmzqtz9XaolMapZ/YZAiQA3p73Ap
PE6u3PzHEORmSCCZ325NpORSPh5/J4uctG0QEKOMrsBf2Xgg/z/vmpi4Mi0aZZPv
3LA1l7ltmI5bQvxvsUM5PaHfLwmESk60t+FL7B9zPTu99YEroCkpPV783BVJJQHV
JHeSycl/uBoBT302VFjLicTTS557B4A11T6zBnTjwiZqeZPkErbZeyt4JNTpAsaz
iTNnuP3DqfD5AF6WRhy5eKw8Kjnm0HIHV+NdYb8dz4XwGgRffZiyjf+6PlNjVJiw
k53FKMcZRwhi2YVReCegDSS+BhxXal0Vrs2rkqbXA2EIMMM//xHjnndcsMP+6MrP
Qtj5NxpQFub0v9JhhNHwxxEofrIYc/ehmS16/BKEe8W5FuX9PMrR/NvGmJNYFvf2
8nz/xMvxoHL7UOHCi/vU4NuDaqsnLEQeha2j6dZm7egso0vYMl7+I5Y1xKpnAZSd
qZH5CI60U3ZuvK89xqOJaqu0czMF4EQc46DpNHYrS7y16pRt1ZiB8UR8AZ1cJHjm
mvPVBuxuQF54PV2Gj478ijI1I+M8jyLul3rgI27/tQiM/2MfeXwg7p7Tgz7sotHG
gChByA4eLk2Xqy+yGvbEttxQ6Zw035dRbvh/6juL8EWchCDFLAPjLwJzt9gwm6tv
1YiqP4uWezHjeItSq+Of/ojcGqLnKqkxUQ/Zmkf/ocSN2VyS47hYgFIt1q/QdJ/V
IMPw2z9uD4cBYGut1MqrIt2dpqfLbXCfihco9M55misuAuejLX5mTwQmzKs3gk+p
gFSy0tnnagMqv2WPolMz8e/eAQDPddCaX0qlkQ8FrmVUK0Qm81mhhO9bKUckmlpm
W1SiQzAfe9A1tTLddS0WckNLD8FsIKaHgcknGg6JVKXjdNR0dG9Y7tY0lxxecC2i
n0q7nsC/Wr3UwTcM3011tz4QPtMzrk5nBTI0gCdEA27MdSOJqvbs9Fp7k9c1GsC3
+O7dANHk5U//wKuqyTNsbiKrAEiyLFRyxK54kPo34sa73WNr925NEcvxKevP8e1s
F1jB6vWGJ+tJLOTOewj+0PzdlHL/lx+fcRA+KrZ8zJClUSPY/uqlt7pujSOKyZaS
xCXNnaW6Zu5WOSQyFCqfcLLLoe1PFmNa25xaRAp67+cuXYJ1tJmtAvS92CrOdDm9
e0k4PP6QEshST0QtrX0X/zbZ0B8/zWDHrF7qhk0+DF4VXCeazE537aXbwoxOZ8Ur
+/JZZsmiti0xH/JsFXXaLcTkbjHQuYGYU2x2B4J3AuQT0uUa7bH4yRvkE56EV7wK
yrStiKIXtQgsevYR+sonbnf/GkqBR8Dy10fs1pr6Y9rB7DmeKqP6Rz865kH8799a
7Cbq9zqS9EgqfOrkNeZCpmuJMhSmVOPPLgRK8+WDFn4X2wM+Shls5XaOgmpJfM6G
UlLyjJnuIYe6Qnr5oXsZanp98RMXN1RQJ4eJLJffh+crLn67PpKd4T61OgoeNN3s
2AsNTqPOEjl9oaddMuxyRGQI9oMn1PUjYoQXmAtSjdoBm4y2M/AWatC7Qy9AEx3c
Ps132KkOtEmqYoA5CN3sdV+G0DHMQGYXy5Xko7jyDDJL8DgFx74CxePYFhdzT9En
/FoiaRVFG3Le749AHr7TmWBHiOO5QnaU33vFhfxwP52FbwnfBOHepmFnmpfEWaOK
I2UpZWnIB3cimPtwyHOmfL2HGLivqpLym8dCvtW+VvRMihI4VGI3nTAYpCcFW07I
A4JRt8+gQNFQUSvJFj3wZcKM8+xPwtSU9LqFLmRwXWX/rHeMvrTMnsbpJTbCa7X/
XvYRH2bkx1EljqvjbWCzMbQ6ZoLumpc+kGUDlWwsdf0bbj8Vd7J9UFJ4hHof+LfW
CXN6FogiD9EPZsuUav+V8s+XIgdAeH2n2DivA8MVbURicdJjFe9536ObkKgFb0w3
pWVY1vVPjb6gtBdpf6KqBrp+9JsNstUkQ99Oyesj8ymotnQv/hB7EqbPCMOJEGCg
DY4ynhhe8nBvIY2kge4KRDB8ispydNqvzoOwVKvP++CfUtEPXpVqEuUHPipPfdnR
zy/u9Rmrz1SnQuABywEqYYODYcVlXXgNmPCFf9Qjyt5bSBKYPH/dwUm0pOIEPQiw
K3CfH8X7GOtMDjgQZGMEar8p1qknrJUDat0WW1QngqRfqDetIZcgxTGQ9d1CXmhZ
cAAtQqlgx3cG+kHAX6ZPwpYtqqDnUMZsJMtguFQMOCb09O40A4IMmzrrnhr0B7bW
J9JP5RARNjhHjhFPrG2WZrdcPGYdUcpakCZBI6hjy+YjIEtKju26AbDMPReQ0OS7
vrGn8AwPJNb3zeJpEi6BOIsbd5BsV1hazsa9JYwS7xHw+ijx9I7SjX9JD5GnuOau
KsRSex21vN1GAnj4+3X5OwX2/FuD/gTt/XPEbay84J3XU34WbimIEVOlQ909zxrd
QncFLXBdlZeQ2spPWKeiFVn7Uhre5kb9lLPpf9Jd2uobQatOYeKGEJxFej6k77uJ
VoZ5MgT5x673LtPMkoxXMVb+sDPXOOnUT6j26yWvcpCkymf4gMN9uezVXd9L1GF/
erwM3blvidYiruDi3gt2qbxqF6g0kR5T2Yd82x70qznyytkKeHPrDvdbaWUOgw2k
j7OVEgFLME/W8QhmmmKP2gws6mHaB8kggCABPu+k5I2OtZ0nltY0K6ORS7GytgJJ
1mKMju2ja1YRh0Mvi7mJottBdY1WWjEiGd6pnDy7HFFSO1SChGxguFKh5XwWfOC4
tjFuHmrabh0kHgt23PrRWV9lD9wfjv9ynxrtGc7kRZU0Agb4a1F/bKmMlAkUf+uj
BwR9uGivRoZJT5n03E4VDG2jSZ5j+E1A/HPcnAFfCnVOeb/2sXAyZtN6fq8+m6ow
Ttj8puqbhhpRRF+mb56Ca8Q7xny4cbDDLZNtghMPuxd6V/bdVXpymDbzYQDvsT9O
n9Gjw+JmbQAt1x5oAbrEtOuhopIB+5+1Lc+WLGGSvGXuJCnH6gjF2oGoTiJkCOgK
augCzpzWcF3w1Dpt7k3HjFoqEXG63HXN7oOummXRH6yqVb6dbO4Lfgp+ZU5EKlox
At2NRFKSPxjJvqvLIUWtT0lbVSPW1Ii3u++CVIBXXZTXyDRR+LHCWnalXyuiN9ek
jaluK13H36pyQv8uxEV5B0EDrdGibQBGs2lbu3XRhfOr1mdDSuZzJ2zQH4Vqs0HT
pf9t/gcGbjX3oDhxif3fzL0wZJz11nBFmNW01QGkYKdJfnmKBl3U5hZ3EwxSJRFm
DTRMlnLCNHj+e5ViKsq1z3/XUdbL2P2np0G70C1rDApcaanSrNiJbsQ11bWNY88d
fByXeW0+0+1ZyCA+WBDhqB5BBvlXKbx+7FjJnF/3Ioa8dobAV8jJDvcNodJZWoYW
00ts0cKUXdHKjsQIcnOPY3CacnwxlevdABwdX6Pp4ReEA1rHYJa0eQ63bHWWVjGi
P5S4pJ6+i09aeKlMQdS/e5Amo/XLCj0UCbj/64JoT3z3HZF/6xj5ohX+K2iDOi/P
uSpqhz/CSF4EfP4UHSZPXXA4vHUjCttXFfERHz0xIu4AqJrDX9FNoXJ+4fr36oYt
HacvPy4zrK7XmZHQNdj4x2FGPdsSv2eWawX145MXBkpLSl9fi4PLUrmtswnba6h3
lUVmxBPVieyGO2c142uEC/lAytiNl+wtcOeOdDkCp1Fk8BlytXxwRdXWA0WLExx6
GBF9EaveNNGk01ewZTawZ2q5ziVtp1FO7nB+WfFekSMBprQ6tekTE+stbP28L5bR
kJMxDLr0kCiB4kiYnoUEiIRUDWUzs0evTBLr3MvC73ZDf7nl+o8xvM3i6Joo2M1D
JfppKKX9a2ITIExffU//aPZ48skt6/FDsGUtRmd+DiHoku7O1TL6wOoU1ITWIYcO
0OE5yIkF2NbtldLIn9t1c8wCVgB9QQ79bBv6J0x/GaNhQ24s4Dr+NwuYLYOQpZlH
n7nxRlebHt7XMSwaiqgN1JyHfit8Up0/Zhpz+Xzfx+76KDzBUbtJIaGuWrWlvZbE
vhz6HgzA1eCiHC1zph+jmbdsIrWle7N37tnIpyS/GPtkWHbX8mB6QbgrMwkVmwLP
6qTfJcf9WJkVBb23Z61b/+sX6lGuqYwaZ823WeheUIr4e6Yqw3QHesBxDNyrgHC2
jCxelkrfHf+X/yXFXzQ/ghtxCzymV3/s5MDETZa/q8l1c3dxl6mWkn6XamY5EevW
sxRKqm8TpKNcDklyBM40hBplps5bsraN+RaD8gCa0GFVUj16izNTCDijFynUyB9L
zqDPoytQq9zUFY97Y51wukTcdgajK+asANOdF1H+uT4k1OJiGo+XpQKNpqfuhZCT
rDxrlog2a83EG+JJK6qKYFQBe+UYOSH34UpjUCp/eLCm1kEGNNhdXsPCkuDv6KMp
5phDy0etDRheMyCZEVBfdrywZJvOmL7r8lJNJPxRU7fciN+xHSrcThiJyPv978B1
Qs+VY1b3lOMbZnTY/yw84IDh9diaLNd5aUmggRh2ZA3x1Q1lbFavTQrGtOvFuFqZ
Wgb6Y+4fne5UbCBqH6Jt2Co2d2C56jygDBAzWmzkmnRlWgSShJy2oQUYVrk4Tmgh
FD5QZtyh7WhAIl3uVEiMNl/6E+j4Kyx6Jgp+FyMAy99UD4LiEy8mcXnPVO7ne1zJ
4D+jbxKLJTE/33bXAyqOVOv/vycWBF876l+khjKutGsY7AjzPHEslAqw+tXPHFAs
6oyYP3WwX0PnSnOK7QQdon7ba9ysNSAsjMDbLpuvsslEx3sanBEZP9niDO+BE+As
lx/YaljxNg7X/9EH9XVpFUDe/MZKrbFHq+Z9vBNkf+gT2h54dI3qm/wbYkllctnu
jGcP7w6k8EeyUc8qfhDoFNkg672EzcGfAuFS3Neby5MhQP2qGLKp78lDEU7zjNh2
OhIpgy/g99qJMOX4/lJJVJIaJz4aMHkPyt0cHrmNuGEqEpppHHdKCWAzVp9NE5Oi
BY21B03yTg99corMFJFU5qTvY0OUMRWoX8OEh5ci8EVSs7HoTuGPEd3ZqdbJ+LLC
U3YyjBORJv0aUotWT0Qocfi+c/9oCZAdyJtSiTiAvLUdAlW4pAMpAW4Co8ckpx9G
N+KaODuK9Hb+PRIHJ0VZATFgxLpswb0MbjoF3EK/FRuDnQONao8p2wKB3nFn68FC
vSh4yFvk0M3wP8kn240/xkEModTXhmhom4Go/9WKHmFZVZYruBgZQpKcrXCZzVR2
j0gPVUxHSMlQ7CkeSjl/Yw9I+OmLdctUengGBUVYqdJ9nZF3lsGVsnlH/xTYkUi6
r8zznz5BEt3/B5CJ8X9Tc/ov/Msvye0QSNBfB8Z6y57rKujjj53ggaSbEPsnH8UJ
reutn/hpgyoKAjqLEJVF+Mg4e69kW6F87vP9dUcPUBkUDvTqLpPhOrVSSExLejA6
usZHNxYwoIKQ0XRv2GO9pqcEVokrYSxsJBSkUdYv/ErQF+Hie3NB0ZwLNO96pmoA
y47aBxQ7LbgNcw5I1YzUiNhG9kvX5BbaqasH0on8xWzMEvTUFjeyajtGpkYFx24a
n/e6weFip0oTivuAe2HK3njn0sgd28hjk5dH6V9Go2gbN1R0g7oWPSPJqd0f3Lvt
b+b9m1zjRr66BYWaWv2Xkw6CRzxGHhYkGwXnuNHY5y+HxCX9szyLUMlJVuBkw+0B
HgSbeprS2VcUZGxJwxI4FP6FbEYALjdZf6mCJTk+99nEwj8JGS8N9ZsfPqUwsX/G
r94wOtli+VZm3am3JVqxZyyaoZNqMP6LOjxrrfFh+Il6bU7GsT1mKNDPP1Wy883s
xXnjSdW1ULzvhdVIvD5JITuc1NjbPFHnas5daTu6PdiE5Y4p4oJxsr36p3Teblx0
oLsHhA2qFC3X29QwadGfU4P/0W8uWCtGJXhKx2q6N5qlCofGQUZPjxZZXqJWpxep
yPL3el26oxA5An1aovsL3s+W8IQeYMqFC/tTLsLF0UErlUyBB1lOCpYq2jsrpDld
CW6rlRW0+Duz4rESOWzlkjeN0Jz+d2eRZUCpDInzDBrTYTd9T95+trp6TSt4Kijp
E8D9nLCQhKIHXl+aUJ9rc2tskOVCITQcHo2kdNbqEfUKj4a4P4SNATUY2U1tWBUI
03mjmMLqvmZZow7o6TxzxK4sfx5TmJsfyUA3m6w3VjXtZbNsgjuIFLjg9Fe9XAku
NRODEiaO5IYNNYyhXfrtsKMGXdwua0DRbH8wfi2U/QPHH4FkvmVJ+9JJNQGOMiiu
cXu8pxaq2cD60HGh3/XhWVUmVKrbtZj1RHKN4RtbdhT8DFhHaapoe0+6DBvIWEd8
/NTkya0Bf9aT9PInE6AB0OpDvsQ6/oLCuxjvpzdF51Low1anP2JluKyXXuV1fn4I
uQNsK4IiOtPjLZ4tEgq6OEo4BydKdkM3Jqn6eBP5ZEQRb2y6/lzS8EKSIQFh9T4Z
BNiqa8buFEzokIFjr9ALp5NkPLvN8c4it1TVB6lvaXp/IEPHndWtzNXcdMoyUVkH
8xgAxcDqR+sildN1Cfy4sGxWaEz66ia5IVCsAUEEmIsVuFnaR/Y3xLB1Ewzl5FTB
rz8Izpzc+AAQ7sbVvwqDuqQkfyr9y69FdBv4uICafyuKTN3pghCX3U83q/0ed8vL
Ng8fifQGe5Dor3dDVjg0yaCsvCStMkJsqc2vZjYPttfHC01rs7pHVyPk4zCCBL0i
c2cKhG8BxLpImMLeYUrWg67hyAvS8TPDFpvGgGRLdxDyc1WVXpT/nLDZxygLnln1
w6FiSh6rf4kWmeg23oxxeP3/H4XZqC3ySHAGMxMeWUybPPMVbCf7gsVloQTJJ2eJ
5hYZaFizwCHu6qVTdJT95Q3emLdmlUripkuG9sMdU9Y1jk9Wj9IGJbRy7nFsemUJ
BcGp/iYFs5i5qHjZVXg1I3GTukI7pn0ZFon6IbYtGSOVR+8gzkQKQZ6aGo6Wj+E/
dIC4JCQ6KSTwnoWd4KgLrXpTtpNBzLIWPcWbcVDPNVWIXogZVXdoCzW/x0a1yNdW
oSMyaNglZtAsWM2HLtgnhdbdPfVhUmGJkj0ePY8hK6a3Ab/tROIPfxjBoi2onujI
rBbKZUUYNg80QJGhWRZAZCGQ2Y5fQw/GSF5ATGFKm1C2q+8A0JHsPGjdheCX9YEh
s30M6EZzs4lc5F+y651qB/BVA2m5T+8M2v7/iCk89BabhbkYUL+rRAd6HcETo0Ik
PexRAZadYTjdKyWO3v4ECx2+AUG8glnrrfRC+DmFwfBeusZHsfOkSA+uhKarhU5a
+T9UgrmwJ1lXc5l26TeZ2RkU1XogBRubNveQwIVj1iwsvQdsDDAznCL8t8AOGW7h
SzVFXv3/Ng85t2tEy8t9vodPsXNIDflTVMrWgmkVhF4q4/SzBL3ii0MD7aY1UNn+
EI31255VfDIjxrgEheSTsdJtEZBU/tScHAT4OWUeolvuHcN33Ac1ov/uoptoVKrn
eqe9F9NPtXoQhoNb2XXhn2NDVahLcJeX4+N+V0X4fW7L55AUJamKzQjGHHmioORc
67ZsSvaKDoW2/wXATq6N3SzIUelSMiWjHNl95YsWhyDlHCH6EE9OpHBuNy8UlH+t
h8ihajHSdEo5vBPaOwtLpRYS2g6BmhKAhyKdM0q7q6NtN1zoT1L7IceMs0FvJ1dI
bhRbTiB2pRk/I0pjIjS4S8gIYSB10z3T2PYRjo16XdQ8z51GSlFl0drbgQdx+Go7
j4AVj8y+xmLmggDBfXqxnLGpnJ1NbylHv1C0AScaW8BLRohhS7GCDpzHpWlcZnkZ
NyQ4G6LOUhD2drOn0pRIbVG5QfELlVuMTivrZiA4PnxGP2I6EzyG1kajvJBS8EVl
XP903AD62khO6exymwA79phM7TwXQPp8Eju5bKG7B9QPI8XAZo3KsvEedgtCJ3Sw
CHAKQNLRy/6+/NmeKmzcktyCo+yl1PSQvEpmWfGEZM/sYx1SxvMNFPrdPk/EFGrL
w9eo70VsXMpKp2NJxQnjpx9lX+Z1iy0FyxlgSCP2IsqMEWFJI8Cu7uanr5wA98KT
JigIXR87AwSfnrfi08eJANVQQLT0hU70L0CJh0zQkIcCgOlJQ1X+FLXH1Bh1iAEy
mFpTTQKfbqeYynZhvmTZN4eHlzXDZ9iUjSjqBCf8maGX3PODl0QiebCO07WUspZm
JA86L5UCKHSz2CPYpGMbGYTdXQIndG+CZZ5R5+XYUGiJRWlsXwGqkIGhhjkBUt92
hSac8V+1P4tn0c32h1rJbBJQXb/vneB++/bsjCoT8BnE0iG5vo+V42pt+18t/dvN
+68UEHT2IhgUjgWcO4eieye5CEcrhwRuwT5rnS8qy+1tinCCCrM8MMx9ZzOCDXC/
3mK1x3raqyD2vPbDjzgIPZxKq5Zwt5gH4lce55gN3cqB2B9XDnZdILd/ipp+0/E7
vBBytdLOZT1K5c//eP/2v1DdWvf5m8tzCkOH8ZnUpMFVVKewbBDn8DyGjiKbb111
fQeMP2pzzRGZvm3zpmXsWTg+qqedUPruU2txGMOVo/BMes7VqsqaUjeAtQaf6dM9
joGrynjWiZSf969XEJUORE7xUM7qRIT+PR3Dl6jJsw9f46rGaI3OYRxsnEcg56j7
t4NpxjiSbw4dK17QDpL9OJXuKrcfROJQCERuw1PLzOz/1vqwFpaMvYjEheyZ3rEK
qyWJUzrRPM7LTnmKMseZ9LxGbO65zw1uKEcRSMOD9LcLURKESRZSdqea8TAfSRGH
IGVS0lM4iHqrXg5DMqIm78sQ/zr08V76KhXvCYPJYCkv9Yz46+D12bqGt5RBELiS
Erzcfbj4Rzts2672KCylf3owqv1nxafgxqXBqeZj1j6ideN6UZc43yBUxr9qlBSk
uGg43fMg0Nts3gLjCnXCeZEEkc1uNSMBSstM2PBUzcYVCY/WUUZVS/OD/UE+2nTZ
4UsGx9geGK56Ir829szCWm+KgudpFkXJiB67/sfqPaVbdB4B2FzI0+EZz7fxoyRZ
FZMBtIyqpIrVo4TY7GFOIinmOuy5c9WXnPlV7xuIYAaNSjLRIX0IU9IGRuuKKKr5
RDxP8pqQmWGVVUUTllqWdeVqFPa3Ajy2AIyOsnnEqvz0jMKIHuGqw3n5oRGhsRV6
evWTcAU6kpRtiK+Ewfxs/0Y+DFl4pNO4p6YHWQaXKoNEg+QBvZAnqGQ6H4hJeME9
VUdK/2sCyJ61XcGcbvzqnI/+O9OjnrTcm48FnHMyK9Lmghsc1kdBEySblMnDfyBK
eFjx+m028jp0Upt/WvPV+qqEAb6OR7vFshyaIdafrTBb2wYaTbTIITGVNZuZhmND
k554MaJDltT8cGytCeck8TWDSOLCwf606Dl0hJIk9L2LomxhPLm/UCM1JyJXQy1N
HX4i+xrm7Oikc3aFcJIkSImwYOPmpo+gobC9w6ogt18v+qARN7PKBOlwQhAU8Xt5
YZwXP3YIJZ/p0Zo7jqY5q188VVJOa8nhra4mMTtm9qz/hiJZfIrmH8iNW1qNakSj
M96fC1YdFbbmvXjGgHf5wIvD04qG++hrefm3CgrxP7eQOz62c/syIuw9Dg3EGEs5
ooU4nXrk7pippKps2o4Oj5WWezcYMIKbNpC4Wb388ylZHRDEhh1ObiluFdCobVCw
IQLWJQKKsmkbC0Y4r/5FJZOqhVCkmYmVGNCmH0PUwBu+6FBj6YMmegQ6w3dIO4JG
62b3AItLCjHr5K9dqanTNa6IvHYLxmO6PQknwLmKvW3Ixsw8IMqkRWdNsSolCDtN
coZJTda7Ue4WJeKkDPBzDc1wVq+hQr60ftAOn7HIaDnLZ9m7halxx04uWQ4BVcdP
zYbTfLI6b/eA4dV8v8mJfFotZhScm/LtVORwNWvMxOsfVqrSAmx2sD7PBG0C5W6q
G6jd8/E1PrNJJvfS64RNKge4Pcexr5BssUiA3czQgKh0n4wS/ZVerthLDZnQQIRX
63Pl1YGpe8PmJYuqkLc0FJrlmjgdTSkhF/7M4WDoo6lxLPQsQmR1WDueTS6yIPeh
kv0npYbIJYhyIjbYSAro41UNTfLSD009fA6TLkKI2N25uuUDL9aXxzZb6QLljLAX
80gD/cn6mfXyDWlAU36+fIqprSqw0uwiswRMrXTANvOp0CFdq454nr1K2AI0xtPS
Rb6cYxlkQnnhskmWaXmx/yABM07DWo+j0ONw3HE1+ALj1fSF/ATLKMKVT+8WNP2T
uQceZ4p47+pudtBG4bk5+fn8fs2CO0jEB62dvtTmrd32zW0Xkarj13m+TF0Satvn
wQO+Kmx8cEWA+DfRkNOEqnsKdqbzuutc+7ZN/jq2Ea7JIIzvWa0Dt0rqJT8igwtP
lsqnTrWgWiAUfmJn8TGdNTRcgVk9L4qXGV3KitDnIF4i8uqBRv6FbTYK8ZEn8IT6
Kzu3ng5+1wuFWTn1srhRAkL75ZZdYnTinZByktRIEefAvGaMzpyuFbzq60hx3XHe
KP0NJuqh/sbv2/FCv97uvH5tGaJQSBJwgeNMypsaKXpexM1EimJwqvBJ7lYCH0WA
8qdrC0IirryOsG1pXeB7QYaWrLy0XaBldTkIQOuQHxrlsp6SaCoZ50EeIifjzeuv
p8mlDKQnty25pwtgRg7zUvdz9V0lqLnNhxW6+Q3MfymiXDzXCxIo4kSHMYA4YrSp
Nft6g0a6TsehVTgpdYQdk3fjgl/Rzp3gbcQVGIP+1P+hdhCQuYH6yP/5XcAnJgzz
q9bPXZnqzJCU8pGLbhWcT8FFZDwXo8rjt7ndcnpkPMiUWg4Y09a9EluMK9UD1HnI
bUZvnz7kJ2SOak9K2BAoSKuVmxod/lJu2dwC7odj/SKczXIN2rJo6w9josnb5o+6
LLALDpFZjiqVLVF50eSAByD+2QlW1KkMRY3fM3+LfL5bHzkk9o3ybsYB19Q4TFzQ
PRw96beo0BR0iqxVfM5SQlc+W7wTTzvumj0Qcc2kkU++3nTDG55wqfliK8BcCMK3
wVCO20XfBdsXHPRHBGFjhM9BLj60cHNUfpM2V2o5z9XYvBqFFXYWTmbQjaTNcO/v
dkAgmUG5WdV48HT6Qrm39AThr/kv/QafISKyguBt6ztCISvo+vspYjp6/0SNE6An
lnD8KPy+FZlK+Kys9/V5PFCDorKqAjmDuzNy0+/kW7IoDUxzs69lYPAggsxwPfOD
m/WhewKw9XsiVam5P88CNhcsagjoIT1P91oIK7x5e/vOh6tImnxm3FefCMvul3MZ
vjo8eSNbF888i7ATaqDBgNcRhT2G8a+kmxi28wmHhy3FwkOdupuHosm7sAFInftQ
m5THBadfeQ6yqF5KfidqlhWF7bgjxoVeLuR0fNUekTMS1k1og14xf7RW3F01CcE1
QG0Oe0yYCuK/Do9MR5yt/tsEPdMHCgi7Zk1lwVh3VdeKV/bkGH3M2OvqGg7czRM2
QPq1DKXPa5jjT2X3PnGT2nw6ZUzilliBsatsBlrvaDuUCXWPvo7QSpgzEkh6X969
9C3w9vLAzKYeb4fsbRRmWFhVgAtVXPxDhP/3LuAZ7LpECJuzxCSpujQYxcZv+9rZ
55INi611cT9aLFC97S0tGL15RmsdLvxWFHp/4jpFMkes9iHs42Rs+K+bo6VqDx8+
pcOaa/B2XnnUrolYN2Op0jvnoe7YcdwN3ozhyiBQkqnjIaApeW58dbvSvTkRTB5/
mvadxuxq4h+UTvPmprh5ojfi+tGgvOkADq+q0Lknd+hYIveHJKd9+0yLQ8dRqjwR
k9Kk4SYcogNDcZIIA8DdNk/s8iClIoUpc4dIiM4GKgkDx1p9oPgGa440EyntZBve
5DNke3986q+Otn3pxp/tpEGziDg0hT4MIz1cvcPsTekmejTVPfvoHPckmUQYkL/P
HlQ7bJZYu1lGYgVGs9V9cH1w+8pOy3QkNKFe8K3T49HUUY2Vc8djyIwrj/XBMhVF
IP/mMzD8advTbrWGxJZzuFN5zskUFOtNpypb0cW3sd+201lG50gAPXkjpHIA5stj
u3q2G7xT9RpOHRAruDSvyBLeDl5jJe/GOF0Azjo+EcrXyPiTFY64h0NvaxpqHmGJ
hIckaCVMDuKd/eZ167mTrnBTcl0wT/MRj41n3mVyNyHpDNEa3ZxWhB59bNSFTjUd
C3iqqmku9sdvOG/U7ESI9j+kUy4WR1MnElW6dYFipXGsxhgUsw4cE8e3GwRVqtc7
f1Pr2dADxzXk48PUfT5/NWGoR7dVoy8CoAQglMT7st5w12HGFhkejnvjiHB30Ggk
V4Fhc1c34lTAzsiZQiRNAzvuBNSF6dzCZqDDUoS34yhmGOPEB0bmc4xhVFh/Hmip
pzirQeSNNXZvNLYDyEJGrcNDst3O707AcfmuKSovy6aPiHRo2c4W1vPRI/P/a2sp
HOF6qD3+iZ6su67R3gcPE/h+W7nRuzi3QYMSB2kTfcznD+AzJx82ennSUlWybKfq
hVkyIoKHO6BoqXCyO9ADW2mQfmdFxiPNnNhnzJcRXhoNvHgsfb5QdYaHwzrrCLxB
axAEjQtIxOPe/G5amK73kZN0hycq7Hw1CUYATl31ax8XLAwz4W4Kxvu/smqHt+WY
FrBUICDFoM9fMrdTRln8BLNp4VeQuJcpJYmKgALIuAIl15AZW7plKfFh4t8850CM
bKHMIDzd2Jwu9+SIT3fUGqvTaqgfUQSkeJCNgNDVIWnIjvpLAAX7thABKxb9c7vZ
zPJg6T+UJ2R0QyVsyiNpU1IKrBnuqzxdH2Y6IdPC1h7MBpynd1wFgEmzZ59iXzGT
onZj6h26KB9SkDrQ6UUYeRPhE8l6leGWPzia+ZvdVgGKE13/rGpBKFTDZz9v7wYz
0LyhjD4QIiRKtH52RGXMONly33GWxNNuQwcLvewl/ka6G+11x7PXMXcurCXdRBds
bW9I04IG6kUWFJ0SUgNknX9T5oWQ32zVK2byRN+hwvOHmEzxp6wbYGr7R1FBGA+S
wMQrSVM9uVGH6wa85RaZ6BUUiNehXPxPkQHQ4Gn5+ezvH3pdPlwoz7laFhXPDFqI
X4NEiuHrLJsJfHJnvwTYqT4dudoocGZmwK6zYUB7DT3Q0jfpNcFQ4mT2F4KMxgm/
fpSdxEE+nCzrRWCNeS3dfdvnrJH04U7x3SaH+x4AfL8RuZOiBHbD32fQ6VPQ6rog
OKLEJjXnhxgKUts/X8nhdtPdnQNV8FDgaGDq9blIPc4Zzg99sn4rLm7EWRt5uS+G
U1KQgQNTj8xbTdhf4ja8/c+dVh4PBaQuSokgO5HMT4OS4lBFgDRcnVRPN2mkz0sW
IIOSeDyXpIWqzrtNSYCkZ6kkAf8fzYD9RXRK+wwF4+h5L7hmvNrbzMAFTK2fHuGx
eLjjo/VVocUo+3L1YMSFv9oU24Cv/vaIfCA10WnJ9iZWoSSdL5zn85fe7br8LZpy
ARpqluur9ZNaYhODcKppSarRAo6fhX3VPSpQRzH0SC1xo/CthZwdUNWaYzu0bN2t
rVsrpcn0ZdcLLgGiDLEP+4Sk6C6sKBNjJY4sukhOpe9Lu68awV7OzBJoglmKNN++
nfQzphE+bWtHSJ/QvsQaRWoMoFaxN/FNhDhE9ZqtvqF/7nobdnEVoY167ETzFAOW
aap3imIZaoAGL9LnOLqvIrTBtL8l2YTJLP3ZkZdlqPa/oNjJW/jkKOdI+S1GSyl9
tvXvOAV8V+jDQPShBwDBUeVFQuNllFR204qTGkjQiglT/QWATRpUe7IjfnnFR8+A
bKTifpVRWX9oeZmYIevjw+RRY2u3JMw2zYZTMAiJKbe2OKyVg8fMRfE4IvR7leeN
BhbMN2R0PMr8y8jlB2BZ6u6snESCi5OoCYQQWoeSNUU4Hv3x3/12+0zkUPKGntKA
vD7XEpg00xBSVFQTQ5r2TF5BG0168Zv+iUIT+46Jpq/XgXV7p8W22WccUpEwxizK
CIioMs3ISCG+GPi17/6LBIUx0PQvLHUDpie6+mZnXp1C7KS7DYKHI9ow/rJ7hk51
xh/+R3YbsDs7RSIfoq9r1XPtIDzYxDyQ4UB5BXQPpWCvDfFRYUqYGqJgDAK0CMh3
CpQlRGXR1sX+zyirUNzzdqvWKdyvyU7DaIu3L0Mu17TH4jyXB1ZTmbjoLjitm2v5
kCup7uKO/C4yb+f0iZxNZOCnMNo6mnI3T15hdjwFyRODOO2TJCGRqJ8iABqL41cd
SdJDeKxthqE7/FMI1u4uTcv8y1hZD1SdF6kn8B9LBNdzkeOdJzWl3/jt11Vsus0m
+BQ81txF/fV6TbUuTS1byQ==
`pragma protect end_protected